--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2018 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--    Generated from core with identifier:                                    --
--    xilinx.com:ip:axi_interconnect:1.06.a                                   --
--                                                                            --
--    The AXI Interconnect core connects one or more AXI4 memory-mapped       --
--    master devices to one AXI4 slave device.                                --
--------------------------------------------------------------------------------
-- Behavioral Simulation Wrapper
-- This file is provided to wrap around the behavioral simulation (if appropriate)

-- Interfaces:
--   AXI4_SLAVE_S00_AXI
--   AXI4_SLAVE_S11_AXI
--   AXI4_SLAVE_S12_AXI
--   AXI4_SLAVE_S10_AXI
--   AXI4_SLAVE_S08_AXI
--   AXI4_SLAVE_S13_AXI
--   AXI4_SLAVE_S02_AXI
--   AXI4_MASTER_M00_AXI
--   AXI4_SLAVE_S15_AXI
--   AXI4_SLAVE_S06_AXI
--   AXI4_SLAVE_S01_AXI
--   AXI4_SLAVE_S09_AXI
--   AXI4_SLAVE_S14_AXI
--   AXI4_SLAVE_S03_AXI
--   AXI4_SLAVE_S04_AXI
--   AXI4_SLAVE_S05_AXI
--   AXI4_SLAVE_S07_AXI

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

LIBRARY axi_interconnect_v1_06_a;
USE axi_interconnect_v1_06_a.axi_interconnect_v1_06_a;

ENTITY axi_fifo_0 IS
  PORT (
    INTERCONNECT_ACLK : IN STD_LOGIC;
    INTERCONNECT_ARESETN : IN STD_LOGIC;
    S00_AXI_ARESET_OUT_N : OUT STD_LOGIC;
    S00_AXI_ACLK : IN STD_LOGIC;
    S00_AXI_AWID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    S00_AXI_AWADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    S00_AXI_AWLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    S00_AXI_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    S00_AXI_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    S00_AXI_AWLOCK : IN STD_LOGIC;
    S00_AXI_AWCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    S00_AXI_AWPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    S00_AXI_AWQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    S00_AXI_AWVALID : IN STD_LOGIC;
    S00_AXI_AWREADY : OUT STD_LOGIC;
    S00_AXI_WDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    S00_AXI_WSTRB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    S00_AXI_WLAST : IN STD_LOGIC;
    S00_AXI_WVALID : IN STD_LOGIC;
    S00_AXI_WREADY : OUT STD_LOGIC;
    S00_AXI_BID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    S00_AXI_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    S00_AXI_BVALID : OUT STD_LOGIC;
    S00_AXI_BREADY : IN STD_LOGIC;
    S00_AXI_ARID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    S00_AXI_ARADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    S00_AXI_ARLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    S00_AXI_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    S00_AXI_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    S00_AXI_ARLOCK : IN STD_LOGIC;
    S00_AXI_ARCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    S00_AXI_ARPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    S00_AXI_ARQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    S00_AXI_ARVALID : IN STD_LOGIC;
    S00_AXI_ARREADY : OUT STD_LOGIC;
    S00_AXI_RID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    S00_AXI_RDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    S00_AXI_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    S00_AXI_RLAST : OUT STD_LOGIC;
    S00_AXI_RVALID : OUT STD_LOGIC;
    S00_AXI_RREADY : IN STD_LOGIC;
    M00_AXI_ARESET_OUT_N : OUT STD_LOGIC;
    M00_AXI_ACLK : IN STD_LOGIC;
    M00_AXI_AWID : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    M00_AXI_AWADDR : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    M00_AXI_AWLEN : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    M00_AXI_AWSIZE : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
    M00_AXI_AWBURST : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    M00_AXI_AWLOCK : OUT STD_LOGIC;
    M00_AXI_AWCACHE : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    M00_AXI_AWPROT : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
    M00_AXI_AWQOS : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    M00_AXI_AWVALID : OUT STD_LOGIC;
    M00_AXI_AWREADY : IN STD_LOGIC;
    M00_AXI_WDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    M00_AXI_WSTRB : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    M00_AXI_WLAST : OUT STD_LOGIC;
    M00_AXI_WVALID : OUT STD_LOGIC;
    M00_AXI_WREADY : IN STD_LOGIC;
    M00_AXI_BID : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    M00_AXI_BRESP : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    M00_AXI_BVALID : IN STD_LOGIC;
    M00_AXI_BREADY : OUT STD_LOGIC;
    M00_AXI_ARID : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    M00_AXI_ARADDR : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    M00_AXI_ARLEN : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    M00_AXI_ARSIZE : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
    M00_AXI_ARBURST : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    M00_AXI_ARLOCK : OUT STD_LOGIC;
    M00_AXI_ARCACHE : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    M00_AXI_ARPROT : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
    M00_AXI_ARQOS : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    M00_AXI_ARVALID : OUT STD_LOGIC;
    M00_AXI_ARREADY : IN STD_LOGIC;
    M00_AXI_RID : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    M00_AXI_RDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    M00_AXI_RRESP : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    M00_AXI_RLAST : IN STD_LOGIC;
    M00_AXI_RVALID : IN STD_LOGIC;
    M00_AXI_RREADY : OUT STD_LOGIC
  );
END axi_fifo_0;

ARCHITECTURE spartan6 OF axi_fifo_0 IS

  constant C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1 : STD_LOGIC_VECTOR(0 DOWNTO 0) := (others => '0');
  constant C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2 : STD_LOGIC_VECTOR(1 DOWNTO 0) := (others => '0');
  constant C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3 : STD_LOGIC_VECTOR(2 DOWNTO 0) := (others => '0');
  constant C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (others => '0');
  constant C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4 : STD_LOGIC_VECTOR(3 DOWNTO 0) := (others => '0');
  constant C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8 : STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '0');

  COMPONENT axi_interconnect_v1_06_a IS
    GENERIC (
      C_FAMILY : STRING;
      C_NUM_SLAVE_PORTS : INTEGER;
      C_THREAD_ID_WIDTH : INTEGER;
      C_THREAD_ID_PORT_WIDTH : INTEGER;
      C_AXI_ADDR_WIDTH : INTEGER;
      C_S00_AXI_DATA_WIDTH : INTEGER;
      C_S01_AXI_DATA_WIDTH : INTEGER;
      C_S02_AXI_DATA_WIDTH : INTEGER;
      C_S03_AXI_DATA_WIDTH : INTEGER;
      C_S04_AXI_DATA_WIDTH : INTEGER;
      C_S05_AXI_DATA_WIDTH : INTEGER;
      C_S06_AXI_DATA_WIDTH : INTEGER;
      C_S07_AXI_DATA_WIDTH : INTEGER;
      C_S08_AXI_DATA_WIDTH : INTEGER;
      C_S09_AXI_DATA_WIDTH : INTEGER;
      C_S10_AXI_DATA_WIDTH : INTEGER;
      C_S11_AXI_DATA_WIDTH : INTEGER;
      C_S12_AXI_DATA_WIDTH : INTEGER;
      C_S13_AXI_DATA_WIDTH : INTEGER;
      C_S14_AXI_DATA_WIDTH : INTEGER;
      C_S15_AXI_DATA_WIDTH : INTEGER;
      C_M00_AXI_DATA_WIDTH : INTEGER;
      C_INTERCONNECT_DATA_WIDTH : INTEGER;
      C_S00_AXI_ACLK_RATIO : STRING;
      C_S01_AXI_ACLK_RATIO : STRING;
      C_S02_AXI_ACLK_RATIO : STRING;
      C_S03_AXI_ACLK_RATIO : STRING;
      C_S04_AXI_ACLK_RATIO : STRING;
      C_S05_AXI_ACLK_RATIO : STRING;
      C_S06_AXI_ACLK_RATIO : STRING;
      C_S07_AXI_ACLK_RATIO : STRING;
      C_S08_AXI_ACLK_RATIO : STRING;
      C_S09_AXI_ACLK_RATIO : STRING;
      C_S10_AXI_ACLK_RATIO : STRING;
      C_S11_AXI_ACLK_RATIO : STRING;
      C_S12_AXI_ACLK_RATIO : STRING;
      C_S13_AXI_ACLK_RATIO : STRING;
      C_S14_AXI_ACLK_RATIO : STRING;
      C_S15_AXI_ACLK_RATIO : STRING;
      C_S00_AXI_IS_ACLK_ASYNC : INTEGER;
      C_S01_AXI_IS_ACLK_ASYNC : INTEGER;
      C_S02_AXI_IS_ACLK_ASYNC : INTEGER;
      C_S03_AXI_IS_ACLK_ASYNC : INTEGER;
      C_S04_AXI_IS_ACLK_ASYNC : INTEGER;
      C_S05_AXI_IS_ACLK_ASYNC : INTEGER;
      C_S06_AXI_IS_ACLK_ASYNC : INTEGER;
      C_S07_AXI_IS_ACLK_ASYNC : INTEGER;
      C_S08_AXI_IS_ACLK_ASYNC : INTEGER;
      C_S09_AXI_IS_ACLK_ASYNC : INTEGER;
      C_S10_AXI_IS_ACLK_ASYNC : INTEGER;
      C_S11_AXI_IS_ACLK_ASYNC : INTEGER;
      C_S12_AXI_IS_ACLK_ASYNC : INTEGER;
      C_S13_AXI_IS_ACLK_ASYNC : INTEGER;
      C_S14_AXI_IS_ACLK_ASYNC : INTEGER;
      C_S15_AXI_IS_ACLK_ASYNC : INTEGER;
      C_M00_AXI_ACLK_RATIO : STRING;
      C_M00_AXI_IS_ACLK_ASYNC : INTEGER;
      C_S00_AXI_READ_WRITE_SUPPORT : STRING;
      C_S01_AXI_READ_WRITE_SUPPORT : STRING;
      C_S02_AXI_READ_WRITE_SUPPORT : STRING;
      C_S03_AXI_READ_WRITE_SUPPORT : STRING;
      C_S04_AXI_READ_WRITE_SUPPORT : STRING;
      C_S05_AXI_READ_WRITE_SUPPORT : STRING;
      C_S06_AXI_READ_WRITE_SUPPORT : STRING;
      C_S07_AXI_READ_WRITE_SUPPORT : STRING;
      C_S08_AXI_READ_WRITE_SUPPORT : STRING;
      C_S09_AXI_READ_WRITE_SUPPORT : STRING;
      C_S10_AXI_READ_WRITE_SUPPORT : STRING;
      C_S11_AXI_READ_WRITE_SUPPORT : STRING;
      C_S12_AXI_READ_WRITE_SUPPORT : STRING;
      C_S13_AXI_READ_WRITE_SUPPORT : STRING;
      C_S14_AXI_READ_WRITE_SUPPORT : STRING;
      C_S15_AXI_READ_WRITE_SUPPORT : STRING;
      C_S00_AXI_WRITE_ACCEPTANCE : INTEGER;
      C_S01_AXI_WRITE_ACCEPTANCE : INTEGER;
      C_S02_AXI_WRITE_ACCEPTANCE : INTEGER;
      C_S03_AXI_WRITE_ACCEPTANCE : INTEGER;
      C_S04_AXI_WRITE_ACCEPTANCE : INTEGER;
      C_S05_AXI_WRITE_ACCEPTANCE : INTEGER;
      C_S06_AXI_WRITE_ACCEPTANCE : INTEGER;
      C_S07_AXI_WRITE_ACCEPTANCE : INTEGER;
      C_S08_AXI_WRITE_ACCEPTANCE : INTEGER;
      C_S09_AXI_WRITE_ACCEPTANCE : INTEGER;
      C_S10_AXI_WRITE_ACCEPTANCE : INTEGER;
      C_S11_AXI_WRITE_ACCEPTANCE : INTEGER;
      C_S12_AXI_WRITE_ACCEPTANCE : INTEGER;
      C_S13_AXI_WRITE_ACCEPTANCE : INTEGER;
      C_S14_AXI_WRITE_ACCEPTANCE : INTEGER;
      C_S15_AXI_WRITE_ACCEPTANCE : INTEGER;
      C_S00_AXI_READ_ACCEPTANCE : INTEGER;
      C_S01_AXI_READ_ACCEPTANCE : INTEGER;
      C_S02_AXI_READ_ACCEPTANCE : INTEGER;
      C_S03_AXI_READ_ACCEPTANCE : INTEGER;
      C_S04_AXI_READ_ACCEPTANCE : INTEGER;
      C_S05_AXI_READ_ACCEPTANCE : INTEGER;
      C_S06_AXI_READ_ACCEPTANCE : INTEGER;
      C_S07_AXI_READ_ACCEPTANCE : INTEGER;
      C_S08_AXI_READ_ACCEPTANCE : INTEGER;
      C_S09_AXI_READ_ACCEPTANCE : INTEGER;
      C_S10_AXI_READ_ACCEPTANCE : INTEGER;
      C_S11_AXI_READ_ACCEPTANCE : INTEGER;
      C_S12_AXI_READ_ACCEPTANCE : INTEGER;
      C_S13_AXI_READ_ACCEPTANCE : INTEGER;
      C_S14_AXI_READ_ACCEPTANCE : INTEGER;
      C_S15_AXI_READ_ACCEPTANCE : INTEGER;
      C_M00_AXI_WRITE_ISSUING : INTEGER;
      C_M00_AXI_READ_ISSUING : INTEGER;
      C_S00_AXI_ARB_PRIORITY : INTEGER;
      C_S01_AXI_ARB_PRIORITY : INTEGER;
      C_S02_AXI_ARB_PRIORITY : INTEGER;
      C_S03_AXI_ARB_PRIORITY : INTEGER;
      C_S04_AXI_ARB_PRIORITY : INTEGER;
      C_S05_AXI_ARB_PRIORITY : INTEGER;
      C_S06_AXI_ARB_PRIORITY : INTEGER;
      C_S07_AXI_ARB_PRIORITY : INTEGER;
      C_S08_AXI_ARB_PRIORITY : INTEGER;
      C_S09_AXI_ARB_PRIORITY : INTEGER;
      C_S10_AXI_ARB_PRIORITY : INTEGER;
      C_S11_AXI_ARB_PRIORITY : INTEGER;
      C_S12_AXI_ARB_PRIORITY : INTEGER;
      C_S13_AXI_ARB_PRIORITY : INTEGER;
      C_S14_AXI_ARB_PRIORITY : INTEGER;
      C_S15_AXI_ARB_PRIORITY : INTEGER;
      C_S00_AXI_WRITE_FIFO_DEPTH : INTEGER;
      C_S01_AXI_WRITE_FIFO_DEPTH : INTEGER;
      C_S02_AXI_WRITE_FIFO_DEPTH : INTEGER;
      C_S03_AXI_WRITE_FIFO_DEPTH : INTEGER;
      C_S04_AXI_WRITE_FIFO_DEPTH : INTEGER;
      C_S05_AXI_WRITE_FIFO_DEPTH : INTEGER;
      C_S06_AXI_WRITE_FIFO_DEPTH : INTEGER;
      C_S07_AXI_WRITE_FIFO_DEPTH : INTEGER;
      C_S08_AXI_WRITE_FIFO_DEPTH : INTEGER;
      C_S09_AXI_WRITE_FIFO_DEPTH : INTEGER;
      C_S10_AXI_WRITE_FIFO_DEPTH : INTEGER;
      C_S11_AXI_WRITE_FIFO_DEPTH : INTEGER;
      C_S12_AXI_WRITE_FIFO_DEPTH : INTEGER;
      C_S13_AXI_WRITE_FIFO_DEPTH : INTEGER;
      C_S14_AXI_WRITE_FIFO_DEPTH : INTEGER;
      C_S15_AXI_WRITE_FIFO_DEPTH : INTEGER;
      C_S00_AXI_READ_FIFO_DEPTH : INTEGER;
      C_S01_AXI_READ_FIFO_DEPTH : INTEGER;
      C_S02_AXI_READ_FIFO_DEPTH : INTEGER;
      C_S03_AXI_READ_FIFO_DEPTH : INTEGER;
      C_S04_AXI_READ_FIFO_DEPTH : INTEGER;
      C_S05_AXI_READ_FIFO_DEPTH : INTEGER;
      C_S06_AXI_READ_FIFO_DEPTH : INTEGER;
      C_S07_AXI_READ_FIFO_DEPTH : INTEGER;
      C_S08_AXI_READ_FIFO_DEPTH : INTEGER;
      C_S09_AXI_READ_FIFO_DEPTH : INTEGER;
      C_S10_AXI_READ_FIFO_DEPTH : INTEGER;
      C_S11_AXI_READ_FIFO_DEPTH : INTEGER;
      C_S12_AXI_READ_FIFO_DEPTH : INTEGER;
      C_S13_AXI_READ_FIFO_DEPTH : INTEGER;
      C_S14_AXI_READ_FIFO_DEPTH : INTEGER;
      C_S15_AXI_READ_FIFO_DEPTH : INTEGER;
      C_M00_AXI_WRITE_FIFO_DEPTH : INTEGER;
      C_M00_AXI_READ_FIFO_DEPTH : INTEGER;
      C_S00_AXI_WRITE_FIFO_DELAY : INTEGER;
      C_S01_AXI_WRITE_FIFO_DELAY : INTEGER;
      C_S02_AXI_WRITE_FIFO_DELAY : INTEGER;
      C_S03_AXI_WRITE_FIFO_DELAY : INTEGER;
      C_S04_AXI_WRITE_FIFO_DELAY : INTEGER;
      C_S05_AXI_WRITE_FIFO_DELAY : INTEGER;
      C_S06_AXI_WRITE_FIFO_DELAY : INTEGER;
      C_S07_AXI_WRITE_FIFO_DELAY : INTEGER;
      C_S08_AXI_WRITE_FIFO_DELAY : INTEGER;
      C_S09_AXI_WRITE_FIFO_DELAY : INTEGER;
      C_S10_AXI_WRITE_FIFO_DELAY : INTEGER;
      C_S11_AXI_WRITE_FIFO_DELAY : INTEGER;
      C_S12_AXI_WRITE_FIFO_DELAY : INTEGER;
      C_S13_AXI_WRITE_FIFO_DELAY : INTEGER;
      C_S14_AXI_WRITE_FIFO_DELAY : INTEGER;
      C_S15_AXI_WRITE_FIFO_DELAY : INTEGER;
      C_S00_AXI_READ_FIFO_DELAY : INTEGER;
      C_S01_AXI_READ_FIFO_DELAY : INTEGER;
      C_S02_AXI_READ_FIFO_DELAY : INTEGER;
      C_S03_AXI_READ_FIFO_DELAY : INTEGER;
      C_S04_AXI_READ_FIFO_DELAY : INTEGER;
      C_S05_AXI_READ_FIFO_DELAY : INTEGER;
      C_S06_AXI_READ_FIFO_DELAY : INTEGER;
      C_S07_AXI_READ_FIFO_DELAY : INTEGER;
      C_S08_AXI_READ_FIFO_DELAY : INTEGER;
      C_S09_AXI_READ_FIFO_DELAY : INTEGER;
      C_S10_AXI_READ_FIFO_DELAY : INTEGER;
      C_S11_AXI_READ_FIFO_DELAY : INTEGER;
      C_S12_AXI_READ_FIFO_DELAY : INTEGER;
      C_S13_AXI_READ_FIFO_DELAY : INTEGER;
      C_S14_AXI_READ_FIFO_DELAY : INTEGER;
      C_S15_AXI_READ_FIFO_DELAY : INTEGER;
      C_M00_AXI_WRITE_FIFO_DELAY : INTEGER;
      C_M00_AXI_READ_FIFO_DELAY : INTEGER;
      C_S00_AXI_REGISTER : INTEGER;
      C_S01_AXI_REGISTER : INTEGER;
      C_S02_AXI_REGISTER : INTEGER;
      C_S03_AXI_REGISTER : INTEGER;
      C_S04_AXI_REGISTER : INTEGER;
      C_S05_AXI_REGISTER : INTEGER;
      C_S06_AXI_REGISTER : INTEGER;
      C_S07_AXI_REGISTER : INTEGER;
      C_S08_AXI_REGISTER : INTEGER;
      C_S09_AXI_REGISTER : INTEGER;
      C_S10_AXI_REGISTER : INTEGER;
      C_S11_AXI_REGISTER : INTEGER;
      C_S12_AXI_REGISTER : INTEGER;
      C_S13_AXI_REGISTER : INTEGER;
      C_S14_AXI_REGISTER : INTEGER;
      C_S15_AXI_REGISTER : INTEGER;
      C_M00_AXI_REGISTER : INTEGER
    );
    PORT (
      INTERCONNECT_ACLK : IN STD_LOGIC;
      INTERCONNECT_ARESETN : IN STD_LOGIC;
      S00_AXI_ARESET_OUT_N : OUT STD_LOGIC;
      S00_AXI_ACLK : IN STD_LOGIC;
      S00_AXI_AWID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S00_AXI_AWADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S00_AXI_AWLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S00_AXI_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S00_AXI_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S00_AXI_AWLOCK : IN STD_LOGIC;
      S00_AXI_AWCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S00_AXI_AWPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S00_AXI_AWQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S00_AXI_AWVALID : IN STD_LOGIC;
      S00_AXI_AWREADY : OUT STD_LOGIC;
      S00_AXI_WDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S00_AXI_WSTRB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S00_AXI_WLAST : IN STD_LOGIC;
      S00_AXI_WVALID : IN STD_LOGIC;
      S00_AXI_WREADY : OUT STD_LOGIC;
      S00_AXI_BID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S00_AXI_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S00_AXI_BVALID : OUT STD_LOGIC;
      S00_AXI_BREADY : IN STD_LOGIC;
      S00_AXI_ARID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S00_AXI_ARADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S00_AXI_ARLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S00_AXI_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S00_AXI_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S00_AXI_ARLOCK : IN STD_LOGIC;
      S00_AXI_ARCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S00_AXI_ARPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S00_AXI_ARQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S00_AXI_ARVALID : IN STD_LOGIC;
      S00_AXI_ARREADY : OUT STD_LOGIC;
      S00_AXI_RID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S00_AXI_RDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      S00_AXI_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S00_AXI_RLAST : OUT STD_LOGIC;
      S00_AXI_RVALID : OUT STD_LOGIC;
      S00_AXI_RREADY : IN STD_LOGIC;
      M00_AXI_ARESET_OUT_N : OUT STD_LOGIC;
      M00_AXI_ACLK : IN STD_LOGIC;
      M00_AXI_AWID : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
      M00_AXI_AWADDR : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      M00_AXI_AWLEN : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
      M00_AXI_AWSIZE : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
      M00_AXI_AWBURST : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      M00_AXI_AWLOCK : OUT STD_LOGIC;
      M00_AXI_AWCACHE : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
      M00_AXI_AWPROT : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
      M00_AXI_AWQOS : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
      M00_AXI_AWVALID : OUT STD_LOGIC;
      M00_AXI_AWREADY : IN STD_LOGIC;
      M00_AXI_WDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      M00_AXI_WSTRB : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
      M00_AXI_WLAST : OUT STD_LOGIC;
      M00_AXI_WVALID : OUT STD_LOGIC;
      M00_AXI_WREADY : IN STD_LOGIC;
      M00_AXI_BID : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      M00_AXI_BRESP : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      M00_AXI_BVALID : IN STD_LOGIC;
      M00_AXI_BREADY : OUT STD_LOGIC;
      M00_AXI_ARID : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
      M00_AXI_ARADDR : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      M00_AXI_ARLEN : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
      M00_AXI_ARSIZE : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
      M00_AXI_ARBURST : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      M00_AXI_ARLOCK : OUT STD_LOGIC;
      M00_AXI_ARCACHE : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
      M00_AXI_ARPROT : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
      M00_AXI_ARQOS : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
      M00_AXI_ARVALID : OUT STD_LOGIC;
      M00_AXI_ARREADY : IN STD_LOGIC;
      M00_AXI_RID : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      M00_AXI_RDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      M00_AXI_RRESP : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      M00_AXI_RLAST : IN STD_LOGIC;
      M00_AXI_RVALID : IN STD_LOGIC;
      M00_AXI_RREADY : OUT STD_LOGIC;
      S01_AXI_ARESET_OUT_N : OUT STD_LOGIC;
      S01_AXI_ACLK : IN STD_LOGIC;
      S01_AXI_AWID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S01_AXI_AWADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S01_AXI_AWLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S01_AXI_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S01_AXI_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S01_AXI_AWLOCK : IN STD_LOGIC;
      S01_AXI_AWCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S01_AXI_AWPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S01_AXI_AWQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S01_AXI_AWVALID : IN STD_LOGIC;
      S01_AXI_AWREADY : OUT STD_LOGIC;
      S01_AXI_WDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S01_AXI_WSTRB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S01_AXI_WLAST : IN STD_LOGIC;
      S01_AXI_WVALID : IN STD_LOGIC;
      S01_AXI_WREADY : OUT STD_LOGIC;
      S01_AXI_BID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S01_AXI_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S01_AXI_BVALID : OUT STD_LOGIC;
      S01_AXI_BREADY : IN STD_LOGIC;
      S01_AXI_ARID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S01_AXI_ARADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S01_AXI_ARLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S01_AXI_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S01_AXI_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S01_AXI_ARLOCK : IN STD_LOGIC;
      S01_AXI_ARCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S01_AXI_ARPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S01_AXI_ARQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S01_AXI_ARVALID : IN STD_LOGIC;
      S01_AXI_ARREADY : OUT STD_LOGIC;
      S01_AXI_RID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S01_AXI_RDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      S01_AXI_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S01_AXI_RLAST : OUT STD_LOGIC;
      S01_AXI_RVALID : OUT STD_LOGIC;
      S01_AXI_RREADY : IN STD_LOGIC;
      S02_AXI_ARESET_OUT_N : OUT STD_LOGIC;
      S02_AXI_ACLK : IN STD_LOGIC;
      S02_AXI_AWID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S02_AXI_AWADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S02_AXI_AWLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S02_AXI_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S02_AXI_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S02_AXI_AWLOCK : IN STD_LOGIC;
      S02_AXI_AWCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S02_AXI_AWPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S02_AXI_AWQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S02_AXI_AWVALID : IN STD_LOGIC;
      S02_AXI_AWREADY : OUT STD_LOGIC;
      S02_AXI_WDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S02_AXI_WSTRB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S02_AXI_WLAST : IN STD_LOGIC;
      S02_AXI_WVALID : IN STD_LOGIC;
      S02_AXI_WREADY : OUT STD_LOGIC;
      S02_AXI_BID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S02_AXI_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S02_AXI_BVALID : OUT STD_LOGIC;
      S02_AXI_BREADY : IN STD_LOGIC;
      S02_AXI_ARID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S02_AXI_ARADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S02_AXI_ARLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S02_AXI_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S02_AXI_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S02_AXI_ARLOCK : IN STD_LOGIC;
      S02_AXI_ARCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S02_AXI_ARPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S02_AXI_ARQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S02_AXI_ARVALID : IN STD_LOGIC;
      S02_AXI_ARREADY : OUT STD_LOGIC;
      S02_AXI_RID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S02_AXI_RDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      S02_AXI_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S02_AXI_RLAST : OUT STD_LOGIC;
      S02_AXI_RVALID : OUT STD_LOGIC;
      S02_AXI_RREADY : IN STD_LOGIC;
      S03_AXI_ARESET_OUT_N : OUT STD_LOGIC;
      S03_AXI_ACLK : IN STD_LOGIC;
      S03_AXI_AWID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S03_AXI_AWADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S03_AXI_AWLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S03_AXI_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S03_AXI_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S03_AXI_AWLOCK : IN STD_LOGIC;
      S03_AXI_AWCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S03_AXI_AWPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S03_AXI_AWQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S03_AXI_AWVALID : IN STD_LOGIC;
      S03_AXI_AWREADY : OUT STD_LOGIC;
      S03_AXI_WDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S03_AXI_WSTRB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S03_AXI_WLAST : IN STD_LOGIC;
      S03_AXI_WVALID : IN STD_LOGIC;
      S03_AXI_WREADY : OUT STD_LOGIC;
      S03_AXI_BID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S03_AXI_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S03_AXI_BVALID : OUT STD_LOGIC;
      S03_AXI_BREADY : IN STD_LOGIC;
      S03_AXI_ARID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S03_AXI_ARADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S03_AXI_ARLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S03_AXI_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S03_AXI_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S03_AXI_ARLOCK : IN STD_LOGIC;
      S03_AXI_ARCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S03_AXI_ARPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S03_AXI_ARQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S03_AXI_ARVALID : IN STD_LOGIC;
      S03_AXI_ARREADY : OUT STD_LOGIC;
      S03_AXI_RID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S03_AXI_RDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      S03_AXI_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S03_AXI_RLAST : OUT STD_LOGIC;
      S03_AXI_RVALID : OUT STD_LOGIC;
      S03_AXI_RREADY : IN STD_LOGIC;
      S04_AXI_ARESET_OUT_N : OUT STD_LOGIC;
      S04_AXI_ACLK : IN STD_LOGIC;
      S04_AXI_AWID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S04_AXI_AWADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S04_AXI_AWLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S04_AXI_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S04_AXI_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S04_AXI_AWLOCK : IN STD_LOGIC;
      S04_AXI_AWCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S04_AXI_AWPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S04_AXI_AWQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S04_AXI_AWVALID : IN STD_LOGIC;
      S04_AXI_AWREADY : OUT STD_LOGIC;
      S04_AXI_WDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S04_AXI_WSTRB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S04_AXI_WLAST : IN STD_LOGIC;
      S04_AXI_WVALID : IN STD_LOGIC;
      S04_AXI_WREADY : OUT STD_LOGIC;
      S04_AXI_BID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S04_AXI_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S04_AXI_BVALID : OUT STD_LOGIC;
      S04_AXI_BREADY : IN STD_LOGIC;
      S04_AXI_ARID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S04_AXI_ARADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S04_AXI_ARLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S04_AXI_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S04_AXI_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S04_AXI_ARLOCK : IN STD_LOGIC;
      S04_AXI_ARCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S04_AXI_ARPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S04_AXI_ARQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S04_AXI_ARVALID : IN STD_LOGIC;
      S04_AXI_ARREADY : OUT STD_LOGIC;
      S04_AXI_RID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S04_AXI_RDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      S04_AXI_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S04_AXI_RLAST : OUT STD_LOGIC;
      S04_AXI_RVALID : OUT STD_LOGIC;
      S04_AXI_RREADY : IN STD_LOGIC;
      S05_AXI_ARESET_OUT_N : OUT STD_LOGIC;
      S05_AXI_ACLK : IN STD_LOGIC;
      S05_AXI_AWID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S05_AXI_AWADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S05_AXI_AWLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S05_AXI_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S05_AXI_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S05_AXI_AWLOCK : IN STD_LOGIC;
      S05_AXI_AWCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S05_AXI_AWPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S05_AXI_AWQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S05_AXI_AWVALID : IN STD_LOGIC;
      S05_AXI_AWREADY : OUT STD_LOGIC;
      S05_AXI_WDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S05_AXI_WSTRB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S05_AXI_WLAST : IN STD_LOGIC;
      S05_AXI_WVALID : IN STD_LOGIC;
      S05_AXI_WREADY : OUT STD_LOGIC;
      S05_AXI_BID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S05_AXI_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S05_AXI_BVALID : OUT STD_LOGIC;
      S05_AXI_BREADY : IN STD_LOGIC;
      S05_AXI_ARID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S05_AXI_ARADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S05_AXI_ARLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S05_AXI_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S05_AXI_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S05_AXI_ARLOCK : IN STD_LOGIC;
      S05_AXI_ARCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S05_AXI_ARPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S05_AXI_ARQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S05_AXI_ARVALID : IN STD_LOGIC;
      S05_AXI_ARREADY : OUT STD_LOGIC;
      S05_AXI_RID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S05_AXI_RDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      S05_AXI_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S05_AXI_RLAST : OUT STD_LOGIC;
      S05_AXI_RVALID : OUT STD_LOGIC;
      S05_AXI_RREADY : IN STD_LOGIC;
      S06_AXI_ARESET_OUT_N : OUT STD_LOGIC;
      S06_AXI_ACLK : IN STD_LOGIC;
      S06_AXI_AWID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S06_AXI_AWADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S06_AXI_AWLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S06_AXI_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S06_AXI_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S06_AXI_AWLOCK : IN STD_LOGIC;
      S06_AXI_AWCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S06_AXI_AWPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S06_AXI_AWQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S06_AXI_AWVALID : IN STD_LOGIC;
      S06_AXI_AWREADY : OUT STD_LOGIC;
      S06_AXI_WDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S06_AXI_WSTRB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S06_AXI_WLAST : IN STD_LOGIC;
      S06_AXI_WVALID : IN STD_LOGIC;
      S06_AXI_WREADY : OUT STD_LOGIC;
      S06_AXI_BID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S06_AXI_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S06_AXI_BVALID : OUT STD_LOGIC;
      S06_AXI_BREADY : IN STD_LOGIC;
      S06_AXI_ARID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S06_AXI_ARADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S06_AXI_ARLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S06_AXI_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S06_AXI_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S06_AXI_ARLOCK : IN STD_LOGIC;
      S06_AXI_ARCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S06_AXI_ARPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S06_AXI_ARQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S06_AXI_ARVALID : IN STD_LOGIC;
      S06_AXI_ARREADY : OUT STD_LOGIC;
      S06_AXI_RID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S06_AXI_RDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      S06_AXI_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S06_AXI_RLAST : OUT STD_LOGIC;
      S06_AXI_RVALID : OUT STD_LOGIC;
      S06_AXI_RREADY : IN STD_LOGIC;
      S07_AXI_ARESET_OUT_N : OUT STD_LOGIC;
      S07_AXI_ACLK : IN STD_LOGIC;
      S07_AXI_AWID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S07_AXI_AWADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S07_AXI_AWLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S07_AXI_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S07_AXI_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S07_AXI_AWLOCK : IN STD_LOGIC;
      S07_AXI_AWCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S07_AXI_AWPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S07_AXI_AWQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S07_AXI_AWVALID : IN STD_LOGIC;
      S07_AXI_AWREADY : OUT STD_LOGIC;
      S07_AXI_WDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S07_AXI_WSTRB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S07_AXI_WLAST : IN STD_LOGIC;
      S07_AXI_WVALID : IN STD_LOGIC;
      S07_AXI_WREADY : OUT STD_LOGIC;
      S07_AXI_BID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S07_AXI_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S07_AXI_BVALID : OUT STD_LOGIC;
      S07_AXI_BREADY : IN STD_LOGIC;
      S07_AXI_ARID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S07_AXI_ARADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S07_AXI_ARLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S07_AXI_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S07_AXI_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S07_AXI_ARLOCK : IN STD_LOGIC;
      S07_AXI_ARCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S07_AXI_ARPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S07_AXI_ARQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S07_AXI_ARVALID : IN STD_LOGIC;
      S07_AXI_ARREADY : OUT STD_LOGIC;
      S07_AXI_RID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S07_AXI_RDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      S07_AXI_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S07_AXI_RLAST : OUT STD_LOGIC;
      S07_AXI_RVALID : OUT STD_LOGIC;
      S07_AXI_RREADY : IN STD_LOGIC;
      S08_AXI_ARESET_OUT_N : OUT STD_LOGIC;
      S08_AXI_ACLK : IN STD_LOGIC;
      S08_AXI_AWID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S08_AXI_AWADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S08_AXI_AWLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S08_AXI_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S08_AXI_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S08_AXI_AWLOCK : IN STD_LOGIC;
      S08_AXI_AWCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S08_AXI_AWPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S08_AXI_AWQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S08_AXI_AWVALID : IN STD_LOGIC;
      S08_AXI_AWREADY : OUT STD_LOGIC;
      S08_AXI_WDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S08_AXI_WSTRB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S08_AXI_WLAST : IN STD_LOGIC;
      S08_AXI_WVALID : IN STD_LOGIC;
      S08_AXI_WREADY : OUT STD_LOGIC;
      S08_AXI_BID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S08_AXI_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S08_AXI_BVALID : OUT STD_LOGIC;
      S08_AXI_BREADY : IN STD_LOGIC;
      S08_AXI_ARID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S08_AXI_ARADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S08_AXI_ARLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S08_AXI_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S08_AXI_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S08_AXI_ARLOCK : IN STD_LOGIC;
      S08_AXI_ARCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S08_AXI_ARPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S08_AXI_ARQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S08_AXI_ARVALID : IN STD_LOGIC;
      S08_AXI_ARREADY : OUT STD_LOGIC;
      S08_AXI_RID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S08_AXI_RDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      S08_AXI_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S08_AXI_RLAST : OUT STD_LOGIC;
      S08_AXI_RVALID : OUT STD_LOGIC;
      S08_AXI_RREADY : IN STD_LOGIC;
      S09_AXI_ARESET_OUT_N : OUT STD_LOGIC;
      S09_AXI_ACLK : IN STD_LOGIC;
      S09_AXI_AWID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S09_AXI_AWADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S09_AXI_AWLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S09_AXI_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S09_AXI_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S09_AXI_AWLOCK : IN STD_LOGIC;
      S09_AXI_AWCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S09_AXI_AWPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S09_AXI_AWQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S09_AXI_AWVALID : IN STD_LOGIC;
      S09_AXI_AWREADY : OUT STD_LOGIC;
      S09_AXI_WDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S09_AXI_WSTRB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S09_AXI_WLAST : IN STD_LOGIC;
      S09_AXI_WVALID : IN STD_LOGIC;
      S09_AXI_WREADY : OUT STD_LOGIC;
      S09_AXI_BID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S09_AXI_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S09_AXI_BVALID : OUT STD_LOGIC;
      S09_AXI_BREADY : IN STD_LOGIC;
      S09_AXI_ARID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S09_AXI_ARADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S09_AXI_ARLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S09_AXI_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S09_AXI_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S09_AXI_ARLOCK : IN STD_LOGIC;
      S09_AXI_ARCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S09_AXI_ARPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S09_AXI_ARQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S09_AXI_ARVALID : IN STD_LOGIC;
      S09_AXI_ARREADY : OUT STD_LOGIC;
      S09_AXI_RID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S09_AXI_RDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      S09_AXI_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S09_AXI_RLAST : OUT STD_LOGIC;
      S09_AXI_RVALID : OUT STD_LOGIC;
      S09_AXI_RREADY : IN STD_LOGIC;
      S10_AXI_ARESET_OUT_N : OUT STD_LOGIC;
      S10_AXI_ACLK : IN STD_LOGIC;
      S10_AXI_AWID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S10_AXI_AWADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S10_AXI_AWLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S10_AXI_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S10_AXI_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S10_AXI_AWLOCK : IN STD_LOGIC;
      S10_AXI_AWCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S10_AXI_AWPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S10_AXI_AWQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S10_AXI_AWVALID : IN STD_LOGIC;
      S10_AXI_AWREADY : OUT STD_LOGIC;
      S10_AXI_WDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S10_AXI_WSTRB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S10_AXI_WLAST : IN STD_LOGIC;
      S10_AXI_WVALID : IN STD_LOGIC;
      S10_AXI_WREADY : OUT STD_LOGIC;
      S10_AXI_BID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S10_AXI_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S10_AXI_BVALID : OUT STD_LOGIC;
      S10_AXI_BREADY : IN STD_LOGIC;
      S10_AXI_ARID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S10_AXI_ARADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S10_AXI_ARLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S10_AXI_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S10_AXI_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S10_AXI_ARLOCK : IN STD_LOGIC;
      S10_AXI_ARCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S10_AXI_ARPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S10_AXI_ARQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S10_AXI_ARVALID : IN STD_LOGIC;
      S10_AXI_ARREADY : OUT STD_LOGIC;
      S10_AXI_RID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S10_AXI_RDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      S10_AXI_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S10_AXI_RLAST : OUT STD_LOGIC;
      S10_AXI_RVALID : OUT STD_LOGIC;
      S10_AXI_RREADY : IN STD_LOGIC;
      S11_AXI_ARESET_OUT_N : OUT STD_LOGIC;
      S11_AXI_ACLK : IN STD_LOGIC;
      S11_AXI_AWID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S11_AXI_AWADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S11_AXI_AWLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S11_AXI_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S11_AXI_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S11_AXI_AWLOCK : IN STD_LOGIC;
      S11_AXI_AWCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S11_AXI_AWPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S11_AXI_AWQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S11_AXI_AWVALID : IN STD_LOGIC;
      S11_AXI_AWREADY : OUT STD_LOGIC;
      S11_AXI_WDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S11_AXI_WSTRB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S11_AXI_WLAST : IN STD_LOGIC;
      S11_AXI_WVALID : IN STD_LOGIC;
      S11_AXI_WREADY : OUT STD_LOGIC;
      S11_AXI_BID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S11_AXI_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S11_AXI_BVALID : OUT STD_LOGIC;
      S11_AXI_BREADY : IN STD_LOGIC;
      S11_AXI_ARID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S11_AXI_ARADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S11_AXI_ARLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S11_AXI_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S11_AXI_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S11_AXI_ARLOCK : IN STD_LOGIC;
      S11_AXI_ARCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S11_AXI_ARPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S11_AXI_ARQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S11_AXI_ARVALID : IN STD_LOGIC;
      S11_AXI_ARREADY : OUT STD_LOGIC;
      S11_AXI_RID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S11_AXI_RDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      S11_AXI_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S11_AXI_RLAST : OUT STD_LOGIC;
      S11_AXI_RVALID : OUT STD_LOGIC;
      S11_AXI_RREADY : IN STD_LOGIC;
      S12_AXI_ARESET_OUT_N : OUT STD_LOGIC;
      S12_AXI_ACLK : IN STD_LOGIC;
      S12_AXI_AWID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S12_AXI_AWADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S12_AXI_AWLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S12_AXI_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S12_AXI_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S12_AXI_AWLOCK : IN STD_LOGIC;
      S12_AXI_AWCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S12_AXI_AWPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S12_AXI_AWQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S12_AXI_AWVALID : IN STD_LOGIC;
      S12_AXI_AWREADY : OUT STD_LOGIC;
      S12_AXI_WDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S12_AXI_WSTRB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S12_AXI_WLAST : IN STD_LOGIC;
      S12_AXI_WVALID : IN STD_LOGIC;
      S12_AXI_WREADY : OUT STD_LOGIC;
      S12_AXI_BID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S12_AXI_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S12_AXI_BVALID : OUT STD_LOGIC;
      S12_AXI_BREADY : IN STD_LOGIC;
      S12_AXI_ARID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S12_AXI_ARADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S12_AXI_ARLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S12_AXI_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S12_AXI_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S12_AXI_ARLOCK : IN STD_LOGIC;
      S12_AXI_ARCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S12_AXI_ARPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S12_AXI_ARQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S12_AXI_ARVALID : IN STD_LOGIC;
      S12_AXI_ARREADY : OUT STD_LOGIC;
      S12_AXI_RID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S12_AXI_RDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      S12_AXI_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S12_AXI_RLAST : OUT STD_LOGIC;
      S12_AXI_RVALID : OUT STD_LOGIC;
      S12_AXI_RREADY : IN STD_LOGIC;
      S13_AXI_ARESET_OUT_N : OUT STD_LOGIC;
      S13_AXI_ACLK : IN STD_LOGIC;
      S13_AXI_AWID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S13_AXI_AWADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S13_AXI_AWLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S13_AXI_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S13_AXI_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S13_AXI_AWLOCK : IN STD_LOGIC;
      S13_AXI_AWCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S13_AXI_AWPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S13_AXI_AWQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S13_AXI_AWVALID : IN STD_LOGIC;
      S13_AXI_AWREADY : OUT STD_LOGIC;
      S13_AXI_WDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S13_AXI_WSTRB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S13_AXI_WLAST : IN STD_LOGIC;
      S13_AXI_WVALID : IN STD_LOGIC;
      S13_AXI_WREADY : OUT STD_LOGIC;
      S13_AXI_BID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S13_AXI_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S13_AXI_BVALID : OUT STD_LOGIC;
      S13_AXI_BREADY : IN STD_LOGIC;
      S13_AXI_ARID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S13_AXI_ARADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S13_AXI_ARLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S13_AXI_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S13_AXI_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S13_AXI_ARLOCK : IN STD_LOGIC;
      S13_AXI_ARCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S13_AXI_ARPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S13_AXI_ARQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S13_AXI_ARVALID : IN STD_LOGIC;
      S13_AXI_ARREADY : OUT STD_LOGIC;
      S13_AXI_RID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S13_AXI_RDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      S13_AXI_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S13_AXI_RLAST : OUT STD_LOGIC;
      S13_AXI_RVALID : OUT STD_LOGIC;
      S13_AXI_RREADY : IN STD_LOGIC;
      S14_AXI_ARESET_OUT_N : OUT STD_LOGIC;
      S14_AXI_ACLK : IN STD_LOGIC;
      S14_AXI_AWID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S14_AXI_AWADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S14_AXI_AWLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S14_AXI_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S14_AXI_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S14_AXI_AWLOCK : IN STD_LOGIC;
      S14_AXI_AWCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S14_AXI_AWPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S14_AXI_AWQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S14_AXI_AWVALID : IN STD_LOGIC;
      S14_AXI_AWREADY : OUT STD_LOGIC;
      S14_AXI_WDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S14_AXI_WSTRB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S14_AXI_WLAST : IN STD_LOGIC;
      S14_AXI_WVALID : IN STD_LOGIC;
      S14_AXI_WREADY : OUT STD_LOGIC;
      S14_AXI_BID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S14_AXI_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S14_AXI_BVALID : OUT STD_LOGIC;
      S14_AXI_BREADY : IN STD_LOGIC;
      S14_AXI_ARID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S14_AXI_ARADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S14_AXI_ARLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S14_AXI_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S14_AXI_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S14_AXI_ARLOCK : IN STD_LOGIC;
      S14_AXI_ARCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S14_AXI_ARPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S14_AXI_ARQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S14_AXI_ARVALID : IN STD_LOGIC;
      S14_AXI_ARREADY : OUT STD_LOGIC;
      S14_AXI_RID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S14_AXI_RDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      S14_AXI_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S14_AXI_RLAST : OUT STD_LOGIC;
      S14_AXI_RVALID : OUT STD_LOGIC;
      S14_AXI_RREADY : IN STD_LOGIC;
      S15_AXI_ARESET_OUT_N : OUT STD_LOGIC;
      S15_AXI_ACLK : IN STD_LOGIC;
      S15_AXI_AWID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S15_AXI_AWADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S15_AXI_AWLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S15_AXI_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S15_AXI_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S15_AXI_AWLOCK : IN STD_LOGIC;
      S15_AXI_AWCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S15_AXI_AWPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S15_AXI_AWQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S15_AXI_AWVALID : IN STD_LOGIC;
      S15_AXI_AWREADY : OUT STD_LOGIC;
      S15_AXI_WDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S15_AXI_WSTRB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S15_AXI_WLAST : IN STD_LOGIC;
      S15_AXI_WVALID : IN STD_LOGIC;
      S15_AXI_WREADY : OUT STD_LOGIC;
      S15_AXI_BID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S15_AXI_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S15_AXI_BVALID : OUT STD_LOGIC;
      S15_AXI_BREADY : IN STD_LOGIC;
      S15_AXI_ARID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S15_AXI_ARADDR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S15_AXI_ARLEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S15_AXI_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S15_AXI_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      S15_AXI_ARLOCK : IN STD_LOGIC;
      S15_AXI_ARCACHE : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S15_AXI_ARPROT : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      S15_AXI_ARQOS : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S15_AXI_ARVALID : IN STD_LOGIC;
      S15_AXI_ARREADY : OUT STD_LOGIC;
      S15_AXI_RID : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      S15_AXI_RDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      S15_AXI_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      S15_AXI_RLAST : OUT STD_LOGIC;
      S15_AXI_RVALID : OUT STD_LOGIC;
      S15_AXI_RREADY : IN STD_LOGIC
    );
  END COMPONENT axi_interconnect_v1_06_a;


  signal DISABLED_OUTPUT_SIGNAL_S01_AXI_ARESET_OUT_N : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S01_AXI_ARREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S01_AXI_AWREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S01_AXI_BID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S01_AXI_BRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S01_AXI_BVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S01_AXI_RDATA : STD_LOGIC_VECTOR(31 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S01_AXI_RID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S01_AXI_RLAST : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S01_AXI_RRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S01_AXI_RVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S01_AXI_WREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S02_AXI_ARESET_OUT_N : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S02_AXI_ARREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S02_AXI_AWREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S02_AXI_BID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S02_AXI_BRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S02_AXI_BVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S02_AXI_RDATA : STD_LOGIC_VECTOR(31 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S02_AXI_RID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S02_AXI_RLAST : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S02_AXI_RRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S02_AXI_RVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S02_AXI_WREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S03_AXI_ARESET_OUT_N : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S03_AXI_ARREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S03_AXI_AWREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S03_AXI_BID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S03_AXI_BRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S03_AXI_BVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S03_AXI_RDATA : STD_LOGIC_VECTOR(31 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S03_AXI_RID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S03_AXI_RLAST : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S03_AXI_RRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S03_AXI_RVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S03_AXI_WREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S04_AXI_ARESET_OUT_N : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S04_AXI_ARREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S04_AXI_AWREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S04_AXI_BID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S04_AXI_BRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S04_AXI_BVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S04_AXI_RDATA : STD_LOGIC_VECTOR(31 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S04_AXI_RID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S04_AXI_RLAST : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S04_AXI_RRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S04_AXI_RVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S04_AXI_WREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S05_AXI_ARESET_OUT_N : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S05_AXI_ARREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S05_AXI_AWREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S05_AXI_BID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S05_AXI_BRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S05_AXI_BVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S05_AXI_RDATA : STD_LOGIC_VECTOR(31 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S05_AXI_RID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S05_AXI_RLAST : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S05_AXI_RRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S05_AXI_RVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S05_AXI_WREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S06_AXI_ARESET_OUT_N : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S06_AXI_ARREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S06_AXI_AWREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S06_AXI_BID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S06_AXI_BRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S06_AXI_BVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S06_AXI_RDATA : STD_LOGIC_VECTOR(31 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S06_AXI_RID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S06_AXI_RLAST : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S06_AXI_RRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S06_AXI_RVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S06_AXI_WREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S07_AXI_ARESET_OUT_N : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S07_AXI_ARREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S07_AXI_AWREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S07_AXI_BID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S07_AXI_BRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S07_AXI_BVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S07_AXI_RDATA : STD_LOGIC_VECTOR(31 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S07_AXI_RID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S07_AXI_RLAST : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S07_AXI_RRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S07_AXI_RVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S07_AXI_WREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S08_AXI_ARESET_OUT_N : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S08_AXI_ARREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S08_AXI_AWREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S08_AXI_BID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S08_AXI_BRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S08_AXI_BVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S08_AXI_RDATA : STD_LOGIC_VECTOR(31 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S08_AXI_RID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S08_AXI_RLAST : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S08_AXI_RRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S08_AXI_RVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S08_AXI_WREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S09_AXI_ARESET_OUT_N : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S09_AXI_ARREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S09_AXI_AWREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S09_AXI_BID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S09_AXI_BRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S09_AXI_BVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S09_AXI_RDATA : STD_LOGIC_VECTOR(31 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S09_AXI_RID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S09_AXI_RLAST : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S09_AXI_RRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S09_AXI_RVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S09_AXI_WREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S10_AXI_ARESET_OUT_N : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S10_AXI_ARREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S10_AXI_AWREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S10_AXI_BID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S10_AXI_BRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S10_AXI_BVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S10_AXI_RDATA : STD_LOGIC_VECTOR(31 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S10_AXI_RID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S10_AXI_RLAST : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S10_AXI_RRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S10_AXI_RVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S10_AXI_WREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S11_AXI_ARESET_OUT_N : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S11_AXI_ARREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S11_AXI_AWREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S11_AXI_BID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S11_AXI_BRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S11_AXI_BVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S11_AXI_RDATA : STD_LOGIC_VECTOR(31 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S11_AXI_RID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S11_AXI_RLAST : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S11_AXI_RRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S11_AXI_RVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S11_AXI_WREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S12_AXI_ARESET_OUT_N : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S12_AXI_ARREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S12_AXI_AWREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S12_AXI_BID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S12_AXI_BRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S12_AXI_BVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S12_AXI_RDATA : STD_LOGIC_VECTOR(31 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S12_AXI_RID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S12_AXI_RLAST : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S12_AXI_RRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S12_AXI_RVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S12_AXI_WREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S13_AXI_ARESET_OUT_N : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S13_AXI_ARREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S13_AXI_AWREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S13_AXI_BID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S13_AXI_BRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S13_AXI_BVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S13_AXI_RDATA : STD_LOGIC_VECTOR(31 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S13_AXI_RID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S13_AXI_RLAST : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S13_AXI_RRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S13_AXI_RVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S13_AXI_WREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S14_AXI_ARESET_OUT_N : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S14_AXI_ARREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S14_AXI_AWREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S14_AXI_BID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S14_AXI_BRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S14_AXI_BVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S14_AXI_RDATA : STD_LOGIC_VECTOR(31 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S14_AXI_RID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S14_AXI_RLAST : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S14_AXI_RRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S14_AXI_RVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S14_AXI_WREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S15_AXI_ARESET_OUT_N : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S15_AXI_ARREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S15_AXI_AWREADY : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S15_AXI_BID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S15_AXI_BRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S15_AXI_BVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S15_AXI_RDATA : STD_LOGIC_VECTOR(31 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S15_AXI_RID : STD_LOGIC_VECTOR(0 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S15_AXI_RLAST : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S15_AXI_RRESP : STD_LOGIC_VECTOR(1 DOWNTO 0);
  signal DISABLED_OUTPUT_SIGNAL_S15_AXI_RVALID : STD_LOGIC;
  signal DISABLED_OUTPUT_SIGNAL_S15_AXI_WREADY : STD_LOGIC;

BEGIN

  U0 : axi_interconnect_v1_06_a
    GENERIC MAP (
      C_AXI_ADDR_WIDTH => 32,
      C_FAMILY => "spartan6",
      C_INTERCONNECT_DATA_WIDTH => 32,
      C_M00_AXI_ACLK_RATIO => "1:1",
      C_M00_AXI_DATA_WIDTH => 32,
      C_M00_AXI_IS_ACLK_ASYNC => 0,
      C_M00_AXI_READ_FIFO_DELAY => 0,
      C_M00_AXI_READ_FIFO_DEPTH => 0,
      C_M00_AXI_READ_ISSUING => 8,
      C_M00_AXI_REGISTER => 0,
      C_M00_AXI_WRITE_FIFO_DELAY => 0,
      C_M00_AXI_WRITE_FIFO_DEPTH => 0,
      C_M00_AXI_WRITE_ISSUING => 8,
      C_NUM_SLAVE_PORTS => 1,
      C_S00_AXI_ACLK_RATIO => "1:1",
      C_S00_AXI_ARB_PRIORITY => 0,
      C_S00_AXI_DATA_WIDTH => 32,
      C_S00_AXI_IS_ACLK_ASYNC => 0,
      C_S00_AXI_READ_ACCEPTANCE => 32,
      C_S00_AXI_READ_FIFO_DELAY => 0,
      C_S00_AXI_READ_FIFO_DEPTH => 0,
      C_S00_AXI_READ_WRITE_SUPPORT => "READ/WRITE",
      C_S00_AXI_REGISTER => 0,
      C_S00_AXI_WRITE_ACCEPTANCE => 32,
      C_S00_AXI_WRITE_FIFO_DELAY => 0,
      C_S00_AXI_WRITE_FIFO_DEPTH => 0,
      C_S01_AXI_ACLK_RATIO => "1:1",
      C_S01_AXI_ARB_PRIORITY => 0,
      C_S01_AXI_DATA_WIDTH => 32,
      C_S01_AXI_IS_ACLK_ASYNC => 0,
      C_S01_AXI_READ_ACCEPTANCE => 1,
      C_S01_AXI_READ_FIFO_DELAY => 0,
      C_S01_AXI_READ_FIFO_DEPTH => 0,
      C_S01_AXI_READ_WRITE_SUPPORT => "READ/WRITE",
      C_S01_AXI_REGISTER => 0,
      C_S01_AXI_WRITE_ACCEPTANCE => 1,
      C_S01_AXI_WRITE_FIFO_DELAY => 0,
      C_S01_AXI_WRITE_FIFO_DEPTH => 0,
      C_S02_AXI_ACLK_RATIO => "1:1",
      C_S02_AXI_ARB_PRIORITY => 0,
      C_S02_AXI_DATA_WIDTH => 32,
      C_S02_AXI_IS_ACLK_ASYNC => 0,
      C_S02_AXI_READ_ACCEPTANCE => 1,
      C_S02_AXI_READ_FIFO_DELAY => 0,
      C_S02_AXI_READ_FIFO_DEPTH => 0,
      C_S02_AXI_READ_WRITE_SUPPORT => "READ/WRITE",
      C_S02_AXI_REGISTER => 0,
      C_S02_AXI_WRITE_ACCEPTANCE => 1,
      C_S02_AXI_WRITE_FIFO_DELAY => 0,
      C_S02_AXI_WRITE_FIFO_DEPTH => 0,
      C_S03_AXI_ACLK_RATIO => "1:1",
      C_S03_AXI_ARB_PRIORITY => 0,
      C_S03_AXI_DATA_WIDTH => 32,
      C_S03_AXI_IS_ACLK_ASYNC => 0,
      C_S03_AXI_READ_ACCEPTANCE => 1,
      C_S03_AXI_READ_FIFO_DELAY => 0,
      C_S03_AXI_READ_FIFO_DEPTH => 0,
      C_S03_AXI_READ_WRITE_SUPPORT => "READ/WRITE",
      C_S03_AXI_REGISTER => 0,
      C_S03_AXI_WRITE_ACCEPTANCE => 1,
      C_S03_AXI_WRITE_FIFO_DELAY => 0,
      C_S03_AXI_WRITE_FIFO_DEPTH => 0,
      C_S04_AXI_ACLK_RATIO => "1:1",
      C_S04_AXI_ARB_PRIORITY => 0,
      C_S04_AXI_DATA_WIDTH => 32,
      C_S04_AXI_IS_ACLK_ASYNC => 0,
      C_S04_AXI_READ_ACCEPTANCE => 1,
      C_S04_AXI_READ_FIFO_DELAY => 0,
      C_S04_AXI_READ_FIFO_DEPTH => 0,
      C_S04_AXI_READ_WRITE_SUPPORT => "READ/WRITE",
      C_S04_AXI_REGISTER => 0,
      C_S04_AXI_WRITE_ACCEPTANCE => 1,
      C_S04_AXI_WRITE_FIFO_DELAY => 0,
      C_S04_AXI_WRITE_FIFO_DEPTH => 0,
      C_S05_AXI_ACLK_RATIO => "1:1",
      C_S05_AXI_ARB_PRIORITY => 0,
      C_S05_AXI_DATA_WIDTH => 32,
      C_S05_AXI_IS_ACLK_ASYNC => 0,
      C_S05_AXI_READ_ACCEPTANCE => 1,
      C_S05_AXI_READ_FIFO_DELAY => 0,
      C_S05_AXI_READ_FIFO_DEPTH => 0,
      C_S05_AXI_READ_WRITE_SUPPORT => "READ/WRITE",
      C_S05_AXI_REGISTER => 0,
      C_S05_AXI_WRITE_ACCEPTANCE => 1,
      C_S05_AXI_WRITE_FIFO_DELAY => 0,
      C_S05_AXI_WRITE_FIFO_DEPTH => 0,
      C_S06_AXI_ACLK_RATIO => "1:1",
      C_S06_AXI_ARB_PRIORITY => 0,
      C_S06_AXI_DATA_WIDTH => 32,
      C_S06_AXI_IS_ACLK_ASYNC => 0,
      C_S06_AXI_READ_ACCEPTANCE => 1,
      C_S06_AXI_READ_FIFO_DELAY => 0,
      C_S06_AXI_READ_FIFO_DEPTH => 0,
      C_S06_AXI_READ_WRITE_SUPPORT => "READ/WRITE",
      C_S06_AXI_REGISTER => 0,
      C_S06_AXI_WRITE_ACCEPTANCE => 1,
      C_S06_AXI_WRITE_FIFO_DELAY => 0,
      C_S06_AXI_WRITE_FIFO_DEPTH => 0,
      C_S07_AXI_ACLK_RATIO => "1:1",
      C_S07_AXI_ARB_PRIORITY => 0,
      C_S07_AXI_DATA_WIDTH => 32,
      C_S07_AXI_IS_ACLK_ASYNC => 0,
      C_S07_AXI_READ_ACCEPTANCE => 1,
      C_S07_AXI_READ_FIFO_DELAY => 0,
      C_S07_AXI_READ_FIFO_DEPTH => 0,
      C_S07_AXI_READ_WRITE_SUPPORT => "READ/WRITE",
      C_S07_AXI_REGISTER => 0,
      C_S07_AXI_WRITE_ACCEPTANCE => 1,
      C_S07_AXI_WRITE_FIFO_DELAY => 0,
      C_S07_AXI_WRITE_FIFO_DEPTH => 0,
      C_S08_AXI_ACLK_RATIO => "1:1",
      C_S08_AXI_ARB_PRIORITY => 0,
      C_S08_AXI_DATA_WIDTH => 32,
      C_S08_AXI_IS_ACLK_ASYNC => 0,
      C_S08_AXI_READ_ACCEPTANCE => 1,
      C_S08_AXI_READ_FIFO_DELAY => 0,
      C_S08_AXI_READ_FIFO_DEPTH => 0,
      C_S08_AXI_READ_WRITE_SUPPORT => "READ/WRITE",
      C_S08_AXI_REGISTER => 0,
      C_S08_AXI_WRITE_ACCEPTANCE => 1,
      C_S08_AXI_WRITE_FIFO_DELAY => 0,
      C_S08_AXI_WRITE_FIFO_DEPTH => 0,
      C_S09_AXI_ACLK_RATIO => "1:1",
      C_S09_AXI_ARB_PRIORITY => 0,
      C_S09_AXI_DATA_WIDTH => 32,
      C_S09_AXI_IS_ACLK_ASYNC => 0,
      C_S09_AXI_READ_ACCEPTANCE => 1,
      C_S09_AXI_READ_FIFO_DELAY => 0,
      C_S09_AXI_READ_FIFO_DEPTH => 0,
      C_S09_AXI_READ_WRITE_SUPPORT => "READ/WRITE",
      C_S09_AXI_REGISTER => 0,
      C_S09_AXI_WRITE_ACCEPTANCE => 1,
      C_S09_AXI_WRITE_FIFO_DELAY => 0,
      C_S09_AXI_WRITE_FIFO_DEPTH => 0,
      C_S10_AXI_ACLK_RATIO => "1:1",
      C_S10_AXI_ARB_PRIORITY => 0,
      C_S10_AXI_DATA_WIDTH => 32,
      C_S10_AXI_IS_ACLK_ASYNC => 0,
      C_S10_AXI_READ_ACCEPTANCE => 1,
      C_S10_AXI_READ_FIFO_DELAY => 0,
      C_S10_AXI_READ_FIFO_DEPTH => 0,
      C_S10_AXI_READ_WRITE_SUPPORT => "READ/WRITE",
      C_S10_AXI_REGISTER => 0,
      C_S10_AXI_WRITE_ACCEPTANCE => 1,
      C_S10_AXI_WRITE_FIFO_DELAY => 0,
      C_S10_AXI_WRITE_FIFO_DEPTH => 0,
      C_S11_AXI_ACLK_RATIO => "1:1",
      C_S11_AXI_ARB_PRIORITY => 0,
      C_S11_AXI_DATA_WIDTH => 32,
      C_S11_AXI_IS_ACLK_ASYNC => 0,
      C_S11_AXI_READ_ACCEPTANCE => 1,
      C_S11_AXI_READ_FIFO_DELAY => 0,
      C_S11_AXI_READ_FIFO_DEPTH => 0,
      C_S11_AXI_READ_WRITE_SUPPORT => "READ/WRITE",
      C_S11_AXI_REGISTER => 0,
      C_S11_AXI_WRITE_ACCEPTANCE => 1,
      C_S11_AXI_WRITE_FIFO_DELAY => 0,
      C_S11_AXI_WRITE_FIFO_DEPTH => 0,
      C_S12_AXI_ACLK_RATIO => "1:1",
      C_S12_AXI_ARB_PRIORITY => 0,
      C_S12_AXI_DATA_WIDTH => 32,
      C_S12_AXI_IS_ACLK_ASYNC => 0,
      C_S12_AXI_READ_ACCEPTANCE => 1,
      C_S12_AXI_READ_FIFO_DELAY => 0,
      C_S12_AXI_READ_FIFO_DEPTH => 0,
      C_S12_AXI_READ_WRITE_SUPPORT => "READ/WRITE",
      C_S12_AXI_REGISTER => 0,
      C_S12_AXI_WRITE_ACCEPTANCE => 1,
      C_S12_AXI_WRITE_FIFO_DELAY => 0,
      C_S12_AXI_WRITE_FIFO_DEPTH => 0,
      C_S13_AXI_ACLK_RATIO => "1:1",
      C_S13_AXI_ARB_PRIORITY => 0,
      C_S13_AXI_DATA_WIDTH => 32,
      C_S13_AXI_IS_ACLK_ASYNC => 0,
      C_S13_AXI_READ_ACCEPTANCE => 1,
      C_S13_AXI_READ_FIFO_DELAY => 0,
      C_S13_AXI_READ_FIFO_DEPTH => 0,
      C_S13_AXI_READ_WRITE_SUPPORT => "READ/WRITE",
      C_S13_AXI_REGISTER => 0,
      C_S13_AXI_WRITE_ACCEPTANCE => 1,
      C_S13_AXI_WRITE_FIFO_DELAY => 0,
      C_S13_AXI_WRITE_FIFO_DEPTH => 0,
      C_S14_AXI_ACLK_RATIO => "1:1",
      C_S14_AXI_ARB_PRIORITY => 0,
      C_S14_AXI_DATA_WIDTH => 32,
      C_S14_AXI_IS_ACLK_ASYNC => 0,
      C_S14_AXI_READ_ACCEPTANCE => 1,
      C_S14_AXI_READ_FIFO_DELAY => 0,
      C_S14_AXI_READ_FIFO_DEPTH => 0,
      C_S14_AXI_READ_WRITE_SUPPORT => "READ/WRITE",
      C_S14_AXI_REGISTER => 0,
      C_S14_AXI_WRITE_ACCEPTANCE => 1,
      C_S14_AXI_WRITE_FIFO_DELAY => 0,
      C_S14_AXI_WRITE_FIFO_DEPTH => 0,
      C_S15_AXI_ACLK_RATIO => "1:1",
      C_S15_AXI_ARB_PRIORITY => 0,
      C_S15_AXI_DATA_WIDTH => 32,
      C_S15_AXI_IS_ACLK_ASYNC => 0,
      C_S15_AXI_READ_ACCEPTANCE => 1,
      C_S15_AXI_READ_FIFO_DELAY => 0,
      C_S15_AXI_READ_FIFO_DEPTH => 0,
      C_S15_AXI_READ_WRITE_SUPPORT => "READ/WRITE",
      C_S15_AXI_REGISTER => 0,
      C_S15_AXI_WRITE_ACCEPTANCE => 1,
      C_S15_AXI_WRITE_FIFO_DELAY => 0,
      C_S15_AXI_WRITE_FIFO_DEPTH => 0,
      C_THREAD_ID_PORT_WIDTH => 1,
      C_THREAD_ID_WIDTH => 0
    )
    PORT MAP (
      INTERCONNECT_ACLK => INTERCONNECT_ACLK,
      INTERCONNECT_ARESETN => INTERCONNECT_ARESETN,
      S00_AXI_ARESET_OUT_N => S00_AXI_ARESET_OUT_N,
      S00_AXI_ACLK => S00_AXI_ACLK,
      S00_AXI_AWID => S00_AXI_AWID,
      S00_AXI_AWADDR => S00_AXI_AWADDR,
      S00_AXI_AWLEN => S00_AXI_AWLEN,
      S00_AXI_AWSIZE => S00_AXI_AWSIZE,
      S00_AXI_AWBURST => S00_AXI_AWBURST,
      S00_AXI_AWLOCK => S00_AXI_AWLOCK,
      S00_AXI_AWCACHE => S00_AXI_AWCACHE,
      S00_AXI_AWPROT => S00_AXI_AWPROT,
      S00_AXI_AWQOS => S00_AXI_AWQOS,
      S00_AXI_AWVALID => S00_AXI_AWVALID,
      S00_AXI_AWREADY => S00_AXI_AWREADY,
      S00_AXI_WDATA => S00_AXI_WDATA,
      S00_AXI_WSTRB => S00_AXI_WSTRB,
      S00_AXI_WLAST => S00_AXI_WLAST,
      S00_AXI_WVALID => S00_AXI_WVALID,
      S00_AXI_WREADY => S00_AXI_WREADY,
      S00_AXI_BID => S00_AXI_BID,
      S00_AXI_BRESP => S00_AXI_BRESP,
      S00_AXI_BVALID => S00_AXI_BVALID,
      S00_AXI_BREADY => S00_AXI_BREADY,
      S00_AXI_ARID => S00_AXI_ARID,
      S00_AXI_ARADDR => S00_AXI_ARADDR,
      S00_AXI_ARLEN => S00_AXI_ARLEN,
      S00_AXI_ARSIZE => S00_AXI_ARSIZE,
      S00_AXI_ARBURST => S00_AXI_ARBURST,
      S00_AXI_ARLOCK => S00_AXI_ARLOCK,
      S00_AXI_ARCACHE => S00_AXI_ARCACHE,
      S00_AXI_ARPROT => S00_AXI_ARPROT,
      S00_AXI_ARQOS => S00_AXI_ARQOS,
      S00_AXI_ARVALID => S00_AXI_ARVALID,
      S00_AXI_ARREADY => S00_AXI_ARREADY,
      S00_AXI_RID => S00_AXI_RID,
      S00_AXI_RDATA => S00_AXI_RDATA,
      S00_AXI_RRESP => S00_AXI_RRESP,
      S00_AXI_RLAST => S00_AXI_RLAST,
      S00_AXI_RVALID => S00_AXI_RVALID,
      S00_AXI_RREADY => S00_AXI_RREADY,
      S01_AXI_ARESET_OUT_N => DISABLED_OUTPUT_SIGNAL_S01_AXI_ARESET_OUT_N,
      S01_AXI_ACLK => '0',
      S01_AXI_AWID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S01_AXI_AWADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S01_AXI_AWLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S01_AXI_AWSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S01_AXI_AWBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S01_AXI_AWLOCK => '0',
      S01_AXI_AWCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S01_AXI_AWPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S01_AXI_AWQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S01_AXI_AWVALID => '0',
      S01_AXI_AWREADY => DISABLED_OUTPUT_SIGNAL_S01_AXI_AWREADY,
      S01_AXI_WDATA => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S01_AXI_WSTRB => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S01_AXI_WLAST => '0',
      S01_AXI_WVALID => '0',
      S01_AXI_WREADY => DISABLED_OUTPUT_SIGNAL_S01_AXI_WREADY,
      S01_AXI_BID => DISABLED_OUTPUT_SIGNAL_S01_AXI_BID,
      S01_AXI_BRESP => DISABLED_OUTPUT_SIGNAL_S01_AXI_BRESP,
      S01_AXI_BVALID => DISABLED_OUTPUT_SIGNAL_S01_AXI_BVALID,
      S01_AXI_BREADY => '0',
      S01_AXI_ARID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S01_AXI_ARADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S01_AXI_ARLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S01_AXI_ARSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S01_AXI_ARBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S01_AXI_ARLOCK => '0',
      S01_AXI_ARCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S01_AXI_ARPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S01_AXI_ARQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S01_AXI_ARVALID => '0',
      S01_AXI_ARREADY => DISABLED_OUTPUT_SIGNAL_S01_AXI_ARREADY,
      S01_AXI_RID => DISABLED_OUTPUT_SIGNAL_S01_AXI_RID,
      S01_AXI_RDATA => DISABLED_OUTPUT_SIGNAL_S01_AXI_RDATA,
      S01_AXI_RRESP => DISABLED_OUTPUT_SIGNAL_S01_AXI_RRESP,
      S01_AXI_RLAST => DISABLED_OUTPUT_SIGNAL_S01_AXI_RLAST,
      S01_AXI_RVALID => DISABLED_OUTPUT_SIGNAL_S01_AXI_RVALID,
      S01_AXI_RREADY => '0',
      S02_AXI_ARESET_OUT_N => DISABLED_OUTPUT_SIGNAL_S02_AXI_ARESET_OUT_N,
      S02_AXI_ACLK => '0',
      S02_AXI_AWID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S02_AXI_AWADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S02_AXI_AWLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S02_AXI_AWSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S02_AXI_AWBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S02_AXI_AWLOCK => '0',
      S02_AXI_AWCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S02_AXI_AWPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S02_AXI_AWQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S02_AXI_AWVALID => '0',
      S02_AXI_AWREADY => DISABLED_OUTPUT_SIGNAL_S02_AXI_AWREADY,
      S02_AXI_WDATA => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S02_AXI_WSTRB => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S02_AXI_WLAST => '0',
      S02_AXI_WVALID => '0',
      S02_AXI_WREADY => DISABLED_OUTPUT_SIGNAL_S02_AXI_WREADY,
      S02_AXI_BID => DISABLED_OUTPUT_SIGNAL_S02_AXI_BID,
      S02_AXI_BRESP => DISABLED_OUTPUT_SIGNAL_S02_AXI_BRESP,
      S02_AXI_BVALID => DISABLED_OUTPUT_SIGNAL_S02_AXI_BVALID,
      S02_AXI_BREADY => '0',
      S02_AXI_ARID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S02_AXI_ARADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S02_AXI_ARLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S02_AXI_ARSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S02_AXI_ARBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S02_AXI_ARLOCK => '0',
      S02_AXI_ARCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S02_AXI_ARPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S02_AXI_ARQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S02_AXI_ARVALID => '0',
      S02_AXI_ARREADY => DISABLED_OUTPUT_SIGNAL_S02_AXI_ARREADY,
      S02_AXI_RID => DISABLED_OUTPUT_SIGNAL_S02_AXI_RID,
      S02_AXI_RDATA => DISABLED_OUTPUT_SIGNAL_S02_AXI_RDATA,
      S02_AXI_RRESP => DISABLED_OUTPUT_SIGNAL_S02_AXI_RRESP,
      S02_AXI_RLAST => DISABLED_OUTPUT_SIGNAL_S02_AXI_RLAST,
      S02_AXI_RVALID => DISABLED_OUTPUT_SIGNAL_S02_AXI_RVALID,
      S02_AXI_RREADY => '0',
      S03_AXI_ARESET_OUT_N => DISABLED_OUTPUT_SIGNAL_S03_AXI_ARESET_OUT_N,
      S03_AXI_ACLK => '0',
      S03_AXI_AWID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S03_AXI_AWADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S03_AXI_AWLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S03_AXI_AWSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S03_AXI_AWBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S03_AXI_AWLOCK => '0',
      S03_AXI_AWCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S03_AXI_AWPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S03_AXI_AWQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S03_AXI_AWVALID => '0',
      S03_AXI_AWREADY => DISABLED_OUTPUT_SIGNAL_S03_AXI_AWREADY,
      S03_AXI_WDATA => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S03_AXI_WSTRB => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S03_AXI_WLAST => '0',
      S03_AXI_WVALID => '0',
      S03_AXI_WREADY => DISABLED_OUTPUT_SIGNAL_S03_AXI_WREADY,
      S03_AXI_BID => DISABLED_OUTPUT_SIGNAL_S03_AXI_BID,
      S03_AXI_BRESP => DISABLED_OUTPUT_SIGNAL_S03_AXI_BRESP,
      S03_AXI_BVALID => DISABLED_OUTPUT_SIGNAL_S03_AXI_BVALID,
      S03_AXI_BREADY => '0',
      S03_AXI_ARID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S03_AXI_ARADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S03_AXI_ARLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S03_AXI_ARSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S03_AXI_ARBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S03_AXI_ARLOCK => '0',
      S03_AXI_ARCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S03_AXI_ARPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S03_AXI_ARQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S03_AXI_ARVALID => '0',
      S03_AXI_ARREADY => DISABLED_OUTPUT_SIGNAL_S03_AXI_ARREADY,
      S03_AXI_RID => DISABLED_OUTPUT_SIGNAL_S03_AXI_RID,
      S03_AXI_RDATA => DISABLED_OUTPUT_SIGNAL_S03_AXI_RDATA,
      S03_AXI_RRESP => DISABLED_OUTPUT_SIGNAL_S03_AXI_RRESP,
      S03_AXI_RLAST => DISABLED_OUTPUT_SIGNAL_S03_AXI_RLAST,
      S03_AXI_RVALID => DISABLED_OUTPUT_SIGNAL_S03_AXI_RVALID,
      S03_AXI_RREADY => '0',
      S04_AXI_ARESET_OUT_N => DISABLED_OUTPUT_SIGNAL_S04_AXI_ARESET_OUT_N,
      S04_AXI_ACLK => '0',
      S04_AXI_AWID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S04_AXI_AWADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S04_AXI_AWLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S04_AXI_AWSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S04_AXI_AWBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S04_AXI_AWLOCK => '0',
      S04_AXI_AWCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S04_AXI_AWPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S04_AXI_AWQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S04_AXI_AWVALID => '0',
      S04_AXI_AWREADY => DISABLED_OUTPUT_SIGNAL_S04_AXI_AWREADY,
      S04_AXI_WDATA => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S04_AXI_WSTRB => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S04_AXI_WLAST => '0',
      S04_AXI_WVALID => '0',
      S04_AXI_WREADY => DISABLED_OUTPUT_SIGNAL_S04_AXI_WREADY,
      S04_AXI_BID => DISABLED_OUTPUT_SIGNAL_S04_AXI_BID,
      S04_AXI_BRESP => DISABLED_OUTPUT_SIGNAL_S04_AXI_BRESP,
      S04_AXI_BVALID => DISABLED_OUTPUT_SIGNAL_S04_AXI_BVALID,
      S04_AXI_BREADY => '0',
      S04_AXI_ARID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S04_AXI_ARADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S04_AXI_ARLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S04_AXI_ARSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S04_AXI_ARBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S04_AXI_ARLOCK => '0',
      S04_AXI_ARCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S04_AXI_ARPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S04_AXI_ARQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S04_AXI_ARVALID => '0',
      S04_AXI_ARREADY => DISABLED_OUTPUT_SIGNAL_S04_AXI_ARREADY,
      S04_AXI_RID => DISABLED_OUTPUT_SIGNAL_S04_AXI_RID,
      S04_AXI_RDATA => DISABLED_OUTPUT_SIGNAL_S04_AXI_RDATA,
      S04_AXI_RRESP => DISABLED_OUTPUT_SIGNAL_S04_AXI_RRESP,
      S04_AXI_RLAST => DISABLED_OUTPUT_SIGNAL_S04_AXI_RLAST,
      S04_AXI_RVALID => DISABLED_OUTPUT_SIGNAL_S04_AXI_RVALID,
      S04_AXI_RREADY => '0',
      S05_AXI_ARESET_OUT_N => DISABLED_OUTPUT_SIGNAL_S05_AXI_ARESET_OUT_N,
      S05_AXI_ACLK => '0',
      S05_AXI_AWID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S05_AXI_AWADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S05_AXI_AWLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S05_AXI_AWSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S05_AXI_AWBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S05_AXI_AWLOCK => '0',
      S05_AXI_AWCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S05_AXI_AWPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S05_AXI_AWQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S05_AXI_AWVALID => '0',
      S05_AXI_AWREADY => DISABLED_OUTPUT_SIGNAL_S05_AXI_AWREADY,
      S05_AXI_WDATA => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S05_AXI_WSTRB => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S05_AXI_WLAST => '0',
      S05_AXI_WVALID => '0',
      S05_AXI_WREADY => DISABLED_OUTPUT_SIGNAL_S05_AXI_WREADY,
      S05_AXI_BID => DISABLED_OUTPUT_SIGNAL_S05_AXI_BID,
      S05_AXI_BRESP => DISABLED_OUTPUT_SIGNAL_S05_AXI_BRESP,
      S05_AXI_BVALID => DISABLED_OUTPUT_SIGNAL_S05_AXI_BVALID,
      S05_AXI_BREADY => '0',
      S05_AXI_ARID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S05_AXI_ARADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S05_AXI_ARLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S05_AXI_ARSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S05_AXI_ARBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S05_AXI_ARLOCK => '0',
      S05_AXI_ARCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S05_AXI_ARPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S05_AXI_ARQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S05_AXI_ARVALID => '0',
      S05_AXI_ARREADY => DISABLED_OUTPUT_SIGNAL_S05_AXI_ARREADY,
      S05_AXI_RID => DISABLED_OUTPUT_SIGNAL_S05_AXI_RID,
      S05_AXI_RDATA => DISABLED_OUTPUT_SIGNAL_S05_AXI_RDATA,
      S05_AXI_RRESP => DISABLED_OUTPUT_SIGNAL_S05_AXI_RRESP,
      S05_AXI_RLAST => DISABLED_OUTPUT_SIGNAL_S05_AXI_RLAST,
      S05_AXI_RVALID => DISABLED_OUTPUT_SIGNAL_S05_AXI_RVALID,
      S05_AXI_RREADY => '0',
      S06_AXI_ARESET_OUT_N => DISABLED_OUTPUT_SIGNAL_S06_AXI_ARESET_OUT_N,
      S06_AXI_ACLK => '0',
      S06_AXI_AWID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S06_AXI_AWADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S06_AXI_AWLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S06_AXI_AWSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S06_AXI_AWBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S06_AXI_AWLOCK => '0',
      S06_AXI_AWCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S06_AXI_AWPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S06_AXI_AWQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S06_AXI_AWVALID => '0',
      S06_AXI_AWREADY => DISABLED_OUTPUT_SIGNAL_S06_AXI_AWREADY,
      S06_AXI_WDATA => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S06_AXI_WSTRB => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S06_AXI_WLAST => '0',
      S06_AXI_WVALID => '0',
      S06_AXI_WREADY => DISABLED_OUTPUT_SIGNAL_S06_AXI_WREADY,
      S06_AXI_BID => DISABLED_OUTPUT_SIGNAL_S06_AXI_BID,
      S06_AXI_BRESP => DISABLED_OUTPUT_SIGNAL_S06_AXI_BRESP,
      S06_AXI_BVALID => DISABLED_OUTPUT_SIGNAL_S06_AXI_BVALID,
      S06_AXI_BREADY => '0',
      S06_AXI_ARID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S06_AXI_ARADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S06_AXI_ARLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S06_AXI_ARSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S06_AXI_ARBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S06_AXI_ARLOCK => '0',
      S06_AXI_ARCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S06_AXI_ARPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S06_AXI_ARQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S06_AXI_ARVALID => '0',
      S06_AXI_ARREADY => DISABLED_OUTPUT_SIGNAL_S06_AXI_ARREADY,
      S06_AXI_RID => DISABLED_OUTPUT_SIGNAL_S06_AXI_RID,
      S06_AXI_RDATA => DISABLED_OUTPUT_SIGNAL_S06_AXI_RDATA,
      S06_AXI_RRESP => DISABLED_OUTPUT_SIGNAL_S06_AXI_RRESP,
      S06_AXI_RLAST => DISABLED_OUTPUT_SIGNAL_S06_AXI_RLAST,
      S06_AXI_RVALID => DISABLED_OUTPUT_SIGNAL_S06_AXI_RVALID,
      S06_AXI_RREADY => '0',
      S07_AXI_ARESET_OUT_N => DISABLED_OUTPUT_SIGNAL_S07_AXI_ARESET_OUT_N,
      S07_AXI_ACLK => '0',
      S07_AXI_AWID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S07_AXI_AWADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S07_AXI_AWLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S07_AXI_AWSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S07_AXI_AWBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S07_AXI_AWLOCK => '0',
      S07_AXI_AWCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S07_AXI_AWPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S07_AXI_AWQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S07_AXI_AWVALID => '0',
      S07_AXI_AWREADY => DISABLED_OUTPUT_SIGNAL_S07_AXI_AWREADY,
      S07_AXI_WDATA => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S07_AXI_WSTRB => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S07_AXI_WLAST => '0',
      S07_AXI_WVALID => '0',
      S07_AXI_WREADY => DISABLED_OUTPUT_SIGNAL_S07_AXI_WREADY,
      S07_AXI_BID => DISABLED_OUTPUT_SIGNAL_S07_AXI_BID,
      S07_AXI_BRESP => DISABLED_OUTPUT_SIGNAL_S07_AXI_BRESP,
      S07_AXI_BVALID => DISABLED_OUTPUT_SIGNAL_S07_AXI_BVALID,
      S07_AXI_BREADY => '0',
      S07_AXI_ARID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S07_AXI_ARADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S07_AXI_ARLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S07_AXI_ARSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S07_AXI_ARBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S07_AXI_ARLOCK => '0',
      S07_AXI_ARCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S07_AXI_ARPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S07_AXI_ARQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S07_AXI_ARVALID => '0',
      S07_AXI_ARREADY => DISABLED_OUTPUT_SIGNAL_S07_AXI_ARREADY,
      S07_AXI_RID => DISABLED_OUTPUT_SIGNAL_S07_AXI_RID,
      S07_AXI_RDATA => DISABLED_OUTPUT_SIGNAL_S07_AXI_RDATA,
      S07_AXI_RRESP => DISABLED_OUTPUT_SIGNAL_S07_AXI_RRESP,
      S07_AXI_RLAST => DISABLED_OUTPUT_SIGNAL_S07_AXI_RLAST,
      S07_AXI_RVALID => DISABLED_OUTPUT_SIGNAL_S07_AXI_RVALID,
      S07_AXI_RREADY => '0',
      S08_AXI_ARESET_OUT_N => DISABLED_OUTPUT_SIGNAL_S08_AXI_ARESET_OUT_N,
      S08_AXI_ACLK => '0',
      S08_AXI_AWID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S08_AXI_AWADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S08_AXI_AWLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S08_AXI_AWSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S08_AXI_AWBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S08_AXI_AWLOCK => '0',
      S08_AXI_AWCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S08_AXI_AWPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S08_AXI_AWQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S08_AXI_AWVALID => '0',
      S08_AXI_AWREADY => DISABLED_OUTPUT_SIGNAL_S08_AXI_AWREADY,
      S08_AXI_WDATA => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S08_AXI_WSTRB => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S08_AXI_WLAST => '0',
      S08_AXI_WVALID => '0',
      S08_AXI_WREADY => DISABLED_OUTPUT_SIGNAL_S08_AXI_WREADY,
      S08_AXI_BID => DISABLED_OUTPUT_SIGNAL_S08_AXI_BID,
      S08_AXI_BRESP => DISABLED_OUTPUT_SIGNAL_S08_AXI_BRESP,
      S08_AXI_BVALID => DISABLED_OUTPUT_SIGNAL_S08_AXI_BVALID,
      S08_AXI_BREADY => '0',
      S08_AXI_ARID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S08_AXI_ARADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S08_AXI_ARLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S08_AXI_ARSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S08_AXI_ARBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S08_AXI_ARLOCK => '0',
      S08_AXI_ARCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S08_AXI_ARPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S08_AXI_ARQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S08_AXI_ARVALID => '0',
      S08_AXI_ARREADY => DISABLED_OUTPUT_SIGNAL_S08_AXI_ARREADY,
      S08_AXI_RID => DISABLED_OUTPUT_SIGNAL_S08_AXI_RID,
      S08_AXI_RDATA => DISABLED_OUTPUT_SIGNAL_S08_AXI_RDATA,
      S08_AXI_RRESP => DISABLED_OUTPUT_SIGNAL_S08_AXI_RRESP,
      S08_AXI_RLAST => DISABLED_OUTPUT_SIGNAL_S08_AXI_RLAST,
      S08_AXI_RVALID => DISABLED_OUTPUT_SIGNAL_S08_AXI_RVALID,
      S08_AXI_RREADY => '0',
      S09_AXI_ARESET_OUT_N => DISABLED_OUTPUT_SIGNAL_S09_AXI_ARESET_OUT_N,
      S09_AXI_ACLK => '0',
      S09_AXI_AWID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S09_AXI_AWADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S09_AXI_AWLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S09_AXI_AWSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S09_AXI_AWBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S09_AXI_AWLOCK => '0',
      S09_AXI_AWCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S09_AXI_AWPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S09_AXI_AWQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S09_AXI_AWVALID => '0',
      S09_AXI_AWREADY => DISABLED_OUTPUT_SIGNAL_S09_AXI_AWREADY,
      S09_AXI_WDATA => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S09_AXI_WSTRB => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S09_AXI_WLAST => '0',
      S09_AXI_WVALID => '0',
      S09_AXI_WREADY => DISABLED_OUTPUT_SIGNAL_S09_AXI_WREADY,
      S09_AXI_BID => DISABLED_OUTPUT_SIGNAL_S09_AXI_BID,
      S09_AXI_BRESP => DISABLED_OUTPUT_SIGNAL_S09_AXI_BRESP,
      S09_AXI_BVALID => DISABLED_OUTPUT_SIGNAL_S09_AXI_BVALID,
      S09_AXI_BREADY => '0',
      S09_AXI_ARID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S09_AXI_ARADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S09_AXI_ARLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S09_AXI_ARSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S09_AXI_ARBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S09_AXI_ARLOCK => '0',
      S09_AXI_ARCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S09_AXI_ARPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S09_AXI_ARQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S09_AXI_ARVALID => '0',
      S09_AXI_ARREADY => DISABLED_OUTPUT_SIGNAL_S09_AXI_ARREADY,
      S09_AXI_RID => DISABLED_OUTPUT_SIGNAL_S09_AXI_RID,
      S09_AXI_RDATA => DISABLED_OUTPUT_SIGNAL_S09_AXI_RDATA,
      S09_AXI_RRESP => DISABLED_OUTPUT_SIGNAL_S09_AXI_RRESP,
      S09_AXI_RLAST => DISABLED_OUTPUT_SIGNAL_S09_AXI_RLAST,
      S09_AXI_RVALID => DISABLED_OUTPUT_SIGNAL_S09_AXI_RVALID,
      S09_AXI_RREADY => '0',
      S10_AXI_ARESET_OUT_N => DISABLED_OUTPUT_SIGNAL_S10_AXI_ARESET_OUT_N,
      S10_AXI_ACLK => '0',
      S10_AXI_AWID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S10_AXI_AWADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S10_AXI_AWLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S10_AXI_AWSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S10_AXI_AWBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S10_AXI_AWLOCK => '0',
      S10_AXI_AWCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S10_AXI_AWPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S10_AXI_AWQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S10_AXI_AWVALID => '0',
      S10_AXI_AWREADY => DISABLED_OUTPUT_SIGNAL_S10_AXI_AWREADY,
      S10_AXI_WDATA => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S10_AXI_WSTRB => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S10_AXI_WLAST => '0',
      S10_AXI_WVALID => '0',
      S10_AXI_WREADY => DISABLED_OUTPUT_SIGNAL_S10_AXI_WREADY,
      S10_AXI_BID => DISABLED_OUTPUT_SIGNAL_S10_AXI_BID,
      S10_AXI_BRESP => DISABLED_OUTPUT_SIGNAL_S10_AXI_BRESP,
      S10_AXI_BVALID => DISABLED_OUTPUT_SIGNAL_S10_AXI_BVALID,
      S10_AXI_BREADY => '0',
      S10_AXI_ARID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S10_AXI_ARADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S10_AXI_ARLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S10_AXI_ARSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S10_AXI_ARBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S10_AXI_ARLOCK => '0',
      S10_AXI_ARCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S10_AXI_ARPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S10_AXI_ARQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S10_AXI_ARVALID => '0',
      S10_AXI_ARREADY => DISABLED_OUTPUT_SIGNAL_S10_AXI_ARREADY,
      S10_AXI_RID => DISABLED_OUTPUT_SIGNAL_S10_AXI_RID,
      S10_AXI_RDATA => DISABLED_OUTPUT_SIGNAL_S10_AXI_RDATA,
      S10_AXI_RRESP => DISABLED_OUTPUT_SIGNAL_S10_AXI_RRESP,
      S10_AXI_RLAST => DISABLED_OUTPUT_SIGNAL_S10_AXI_RLAST,
      S10_AXI_RVALID => DISABLED_OUTPUT_SIGNAL_S10_AXI_RVALID,
      S10_AXI_RREADY => '0',
      S11_AXI_ARESET_OUT_N => DISABLED_OUTPUT_SIGNAL_S11_AXI_ARESET_OUT_N,
      S11_AXI_ACLK => '0',
      S11_AXI_AWID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S11_AXI_AWADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S11_AXI_AWLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S11_AXI_AWSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S11_AXI_AWBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S11_AXI_AWLOCK => '0',
      S11_AXI_AWCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S11_AXI_AWPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S11_AXI_AWQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S11_AXI_AWVALID => '0',
      S11_AXI_AWREADY => DISABLED_OUTPUT_SIGNAL_S11_AXI_AWREADY,
      S11_AXI_WDATA => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S11_AXI_WSTRB => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S11_AXI_WLAST => '0',
      S11_AXI_WVALID => '0',
      S11_AXI_WREADY => DISABLED_OUTPUT_SIGNAL_S11_AXI_WREADY,
      S11_AXI_BID => DISABLED_OUTPUT_SIGNAL_S11_AXI_BID,
      S11_AXI_BRESP => DISABLED_OUTPUT_SIGNAL_S11_AXI_BRESP,
      S11_AXI_BVALID => DISABLED_OUTPUT_SIGNAL_S11_AXI_BVALID,
      S11_AXI_BREADY => '0',
      S11_AXI_ARID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S11_AXI_ARADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S11_AXI_ARLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S11_AXI_ARSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S11_AXI_ARBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S11_AXI_ARLOCK => '0',
      S11_AXI_ARCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S11_AXI_ARPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S11_AXI_ARQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S11_AXI_ARVALID => '0',
      S11_AXI_ARREADY => DISABLED_OUTPUT_SIGNAL_S11_AXI_ARREADY,
      S11_AXI_RID => DISABLED_OUTPUT_SIGNAL_S11_AXI_RID,
      S11_AXI_RDATA => DISABLED_OUTPUT_SIGNAL_S11_AXI_RDATA,
      S11_AXI_RRESP => DISABLED_OUTPUT_SIGNAL_S11_AXI_RRESP,
      S11_AXI_RLAST => DISABLED_OUTPUT_SIGNAL_S11_AXI_RLAST,
      S11_AXI_RVALID => DISABLED_OUTPUT_SIGNAL_S11_AXI_RVALID,
      S11_AXI_RREADY => '0',
      S12_AXI_ARESET_OUT_N => DISABLED_OUTPUT_SIGNAL_S12_AXI_ARESET_OUT_N,
      S12_AXI_ACLK => '0',
      S12_AXI_AWID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S12_AXI_AWADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S12_AXI_AWLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S12_AXI_AWSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S12_AXI_AWBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S12_AXI_AWLOCK => '0',
      S12_AXI_AWCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S12_AXI_AWPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S12_AXI_AWQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S12_AXI_AWVALID => '0',
      S12_AXI_AWREADY => DISABLED_OUTPUT_SIGNAL_S12_AXI_AWREADY,
      S12_AXI_WDATA => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S12_AXI_WSTRB => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S12_AXI_WLAST => '0',
      S12_AXI_WVALID => '0',
      S12_AXI_WREADY => DISABLED_OUTPUT_SIGNAL_S12_AXI_WREADY,
      S12_AXI_BID => DISABLED_OUTPUT_SIGNAL_S12_AXI_BID,
      S12_AXI_BRESP => DISABLED_OUTPUT_SIGNAL_S12_AXI_BRESP,
      S12_AXI_BVALID => DISABLED_OUTPUT_SIGNAL_S12_AXI_BVALID,
      S12_AXI_BREADY => '0',
      S12_AXI_ARID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S12_AXI_ARADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S12_AXI_ARLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S12_AXI_ARSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S12_AXI_ARBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S12_AXI_ARLOCK => '0',
      S12_AXI_ARCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S12_AXI_ARPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S12_AXI_ARQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S12_AXI_ARVALID => '0',
      S12_AXI_ARREADY => DISABLED_OUTPUT_SIGNAL_S12_AXI_ARREADY,
      S12_AXI_RID => DISABLED_OUTPUT_SIGNAL_S12_AXI_RID,
      S12_AXI_RDATA => DISABLED_OUTPUT_SIGNAL_S12_AXI_RDATA,
      S12_AXI_RRESP => DISABLED_OUTPUT_SIGNAL_S12_AXI_RRESP,
      S12_AXI_RLAST => DISABLED_OUTPUT_SIGNAL_S12_AXI_RLAST,
      S12_AXI_RVALID => DISABLED_OUTPUT_SIGNAL_S12_AXI_RVALID,
      S12_AXI_RREADY => '0',
      S13_AXI_ARESET_OUT_N => DISABLED_OUTPUT_SIGNAL_S13_AXI_ARESET_OUT_N,
      S13_AXI_ACLK => '0',
      S13_AXI_AWID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S13_AXI_AWADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S13_AXI_AWLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S13_AXI_AWSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S13_AXI_AWBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S13_AXI_AWLOCK => '0',
      S13_AXI_AWCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S13_AXI_AWPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S13_AXI_AWQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S13_AXI_AWVALID => '0',
      S13_AXI_AWREADY => DISABLED_OUTPUT_SIGNAL_S13_AXI_AWREADY,
      S13_AXI_WDATA => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S13_AXI_WSTRB => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S13_AXI_WLAST => '0',
      S13_AXI_WVALID => '0',
      S13_AXI_WREADY => DISABLED_OUTPUT_SIGNAL_S13_AXI_WREADY,
      S13_AXI_BID => DISABLED_OUTPUT_SIGNAL_S13_AXI_BID,
      S13_AXI_BRESP => DISABLED_OUTPUT_SIGNAL_S13_AXI_BRESP,
      S13_AXI_BVALID => DISABLED_OUTPUT_SIGNAL_S13_AXI_BVALID,
      S13_AXI_BREADY => '0',
      S13_AXI_ARID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S13_AXI_ARADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S13_AXI_ARLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S13_AXI_ARSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S13_AXI_ARBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S13_AXI_ARLOCK => '0',
      S13_AXI_ARCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S13_AXI_ARPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S13_AXI_ARQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S13_AXI_ARVALID => '0',
      S13_AXI_ARREADY => DISABLED_OUTPUT_SIGNAL_S13_AXI_ARREADY,
      S13_AXI_RID => DISABLED_OUTPUT_SIGNAL_S13_AXI_RID,
      S13_AXI_RDATA => DISABLED_OUTPUT_SIGNAL_S13_AXI_RDATA,
      S13_AXI_RRESP => DISABLED_OUTPUT_SIGNAL_S13_AXI_RRESP,
      S13_AXI_RLAST => DISABLED_OUTPUT_SIGNAL_S13_AXI_RLAST,
      S13_AXI_RVALID => DISABLED_OUTPUT_SIGNAL_S13_AXI_RVALID,
      S13_AXI_RREADY => '0',
      S14_AXI_ARESET_OUT_N => DISABLED_OUTPUT_SIGNAL_S14_AXI_ARESET_OUT_N,
      S14_AXI_ACLK => '0',
      S14_AXI_AWID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S14_AXI_AWADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S14_AXI_AWLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S14_AXI_AWSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S14_AXI_AWBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S14_AXI_AWLOCK => '0',
      S14_AXI_AWCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S14_AXI_AWPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S14_AXI_AWQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S14_AXI_AWVALID => '0',
      S14_AXI_AWREADY => DISABLED_OUTPUT_SIGNAL_S14_AXI_AWREADY,
      S14_AXI_WDATA => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S14_AXI_WSTRB => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S14_AXI_WLAST => '0',
      S14_AXI_WVALID => '0',
      S14_AXI_WREADY => DISABLED_OUTPUT_SIGNAL_S14_AXI_WREADY,
      S14_AXI_BID => DISABLED_OUTPUT_SIGNAL_S14_AXI_BID,
      S14_AXI_BRESP => DISABLED_OUTPUT_SIGNAL_S14_AXI_BRESP,
      S14_AXI_BVALID => DISABLED_OUTPUT_SIGNAL_S14_AXI_BVALID,
      S14_AXI_BREADY => '0',
      S14_AXI_ARID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S14_AXI_ARADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S14_AXI_ARLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S14_AXI_ARSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S14_AXI_ARBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S14_AXI_ARLOCK => '0',
      S14_AXI_ARCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S14_AXI_ARPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S14_AXI_ARQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S14_AXI_ARVALID => '0',
      S14_AXI_ARREADY => DISABLED_OUTPUT_SIGNAL_S14_AXI_ARREADY,
      S14_AXI_RID => DISABLED_OUTPUT_SIGNAL_S14_AXI_RID,
      S14_AXI_RDATA => DISABLED_OUTPUT_SIGNAL_S14_AXI_RDATA,
      S14_AXI_RRESP => DISABLED_OUTPUT_SIGNAL_S14_AXI_RRESP,
      S14_AXI_RLAST => DISABLED_OUTPUT_SIGNAL_S14_AXI_RLAST,
      S14_AXI_RVALID => DISABLED_OUTPUT_SIGNAL_S14_AXI_RVALID,
      S14_AXI_RREADY => '0',
      S15_AXI_ARESET_OUT_N => DISABLED_OUTPUT_SIGNAL_S15_AXI_ARESET_OUT_N,
      S15_AXI_ACLK => '0',
      S15_AXI_AWID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S15_AXI_AWADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S15_AXI_AWLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S15_AXI_AWSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S15_AXI_AWBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S15_AXI_AWLOCK => '0',
      S15_AXI_AWCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S15_AXI_AWPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S15_AXI_AWQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S15_AXI_AWVALID => '0',
      S15_AXI_AWREADY => DISABLED_OUTPUT_SIGNAL_S15_AXI_AWREADY,
      S15_AXI_WDATA => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S15_AXI_WSTRB => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S15_AXI_WLAST => '0',
      S15_AXI_WVALID => '0',
      S15_AXI_WREADY => DISABLED_OUTPUT_SIGNAL_S15_AXI_WREADY,
      S15_AXI_BID => DISABLED_OUTPUT_SIGNAL_S15_AXI_BID,
      S15_AXI_BRESP => DISABLED_OUTPUT_SIGNAL_S15_AXI_BRESP,
      S15_AXI_BVALID => DISABLED_OUTPUT_SIGNAL_S15_AXI_BVALID,
      S15_AXI_BREADY => '0',
      S15_AXI_ARID => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_1,
      S15_AXI_ARADDR => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_32,
      S15_AXI_ARLEN => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_8,
      S15_AXI_ARSIZE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S15_AXI_ARBURST => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_2,
      S15_AXI_ARLOCK => '0',
      S15_AXI_ARCACHE => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S15_AXI_ARPROT => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_3,
      S15_AXI_ARQOS => C_DEFAULT_INPUT_DRIVER_AGGREGATION_SIGNAL_4,
      S15_AXI_ARVALID => '0',
      S15_AXI_ARREADY => DISABLED_OUTPUT_SIGNAL_S15_AXI_ARREADY,
      S15_AXI_RID => DISABLED_OUTPUT_SIGNAL_S15_AXI_RID,
      S15_AXI_RDATA => DISABLED_OUTPUT_SIGNAL_S15_AXI_RDATA,
      S15_AXI_RRESP => DISABLED_OUTPUT_SIGNAL_S15_AXI_RRESP,
      S15_AXI_RLAST => DISABLED_OUTPUT_SIGNAL_S15_AXI_RLAST,
      S15_AXI_RVALID => DISABLED_OUTPUT_SIGNAL_S15_AXI_RVALID,
      S15_AXI_RREADY => '0',
      M00_AXI_ARESET_OUT_N => M00_AXI_ARESET_OUT_N,
      M00_AXI_ACLK => M00_AXI_ACLK,
      M00_AXI_AWID => M00_AXI_AWID,
      M00_AXI_AWADDR => M00_AXI_AWADDR,
      M00_AXI_AWLEN => M00_AXI_AWLEN,
      M00_AXI_AWSIZE => M00_AXI_AWSIZE,
      M00_AXI_AWBURST => M00_AXI_AWBURST,
      M00_AXI_AWLOCK => M00_AXI_AWLOCK,
      M00_AXI_AWCACHE => M00_AXI_AWCACHE,
      M00_AXI_AWPROT => M00_AXI_AWPROT,
      M00_AXI_AWQOS => M00_AXI_AWQOS,
      M00_AXI_AWVALID => M00_AXI_AWVALID,
      M00_AXI_AWREADY => M00_AXI_AWREADY,
      M00_AXI_WDATA => M00_AXI_WDATA,
      M00_AXI_WSTRB => M00_AXI_WSTRB,
      M00_AXI_WLAST => M00_AXI_WLAST,
      M00_AXI_WVALID => M00_AXI_WVALID,
      M00_AXI_WREADY => M00_AXI_WREADY,
      M00_AXI_BID => M00_AXI_BID,
      M00_AXI_BRESP => M00_AXI_BRESP,
      M00_AXI_BVALID => M00_AXI_BVALID,
      M00_AXI_BREADY => M00_AXI_BREADY,
      M00_AXI_ARID => M00_AXI_ARID,
      M00_AXI_ARADDR => M00_AXI_ARADDR,
      M00_AXI_ARLEN => M00_AXI_ARLEN,
      M00_AXI_ARSIZE => M00_AXI_ARSIZE,
      M00_AXI_ARBURST => M00_AXI_ARBURST,
      M00_AXI_ARLOCK => M00_AXI_ARLOCK,
      M00_AXI_ARCACHE => M00_AXI_ARCACHE,
      M00_AXI_ARPROT => M00_AXI_ARPROT,
      M00_AXI_ARQOS => M00_AXI_ARQOS,
      M00_AXI_ARVALID => M00_AXI_ARVALID,
      M00_AXI_ARREADY => M00_AXI_ARREADY,
      M00_AXI_RID => M00_AXI_RID,
      M00_AXI_RDATA => M00_AXI_RDATA,
      M00_AXI_RRESP => M00_AXI_RRESP,
      M00_AXI_RLAST => M00_AXI_RLAST,
      M00_AXI_RVALID => M00_AXI_RVALID,
      M00_AXI_RREADY => M00_AXI_RREADY
    );

END spartan6;
