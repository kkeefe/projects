--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2018 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--    Generated from core with identifier:                                    --
--    xilinx.com:ip:axis_interconnect:1.1                                     --
--                                                                            --
--    The AXI4-Stream Interconnect IP provides the infrastructure to          --
--    connect multiple AXI4-Stream masters and slaves.  The configurable      --
--    interconnect features a 16x16 switch, data FIFOs, register slices,      --
--    data width converters and clock rate converters.                        --
--------------------------------------------------------------------------------
-- Source Code Wrapper
-- This file is provided to wrap around the source code (if appropriate)

-- Interfaces:
--   S00_AXIS
--   S01_AXIS
--   S02_AXIS
--   S03_AXIS
--   S04_AXIS
--   S05_AXIS
--   S06_AXIS
--   S07_AXIS
--   S08_AXIS
--   S09_AXIS
--   S10_AXIS
--   S11_AXIS
--   S12_AXIS
--   S13_AXIS
--   S14_AXIS
--   S15_AXIS
--   M00_AXIS
--   M01_AXIS
--   M02_AXIS
--   M03_AXIS
--   M04_AXIS
--   M05_AXIS
--   M06_AXIS
--   M07_AXIS
--   M08_AXIS
--   M09_AXIS
--   M10_AXIS
--   M11_AXIS
--   M12_AXIS
--   M13_AXIS
--   M14_AXIS
--   M15_AXIS
--   RSTIF
--   CLKIF
--   CLKENIF
--   S00_RSTIF
--   S00_CLKIF
--   S00_CLKENIF
--   M00_RSTIF
--   M00_CLKIF
--   M00_CLKENIF
--   S01_RSTIF
--   S01_CLKIF
--   S01_CLKENIF
--   M01_RSTIF
--   M01_CLKIF
--   M01_CLKENIF
--   S02_RSTIF
--   S02_CLKIF
--   S02_CLKENIF
--   M02_RSTIF
--   M02_CLKIF
--   M02_CLKENIF
--   S03_RSTIF
--   S03_CLKIF
--   S03_CLKENIF
--   M03_RSTIF
--   M03_CLKIF
--   M03_CLKENIF
--   S04_RSTIF
--   S04_CLKIF
--   S04_CLKENIF
--   M04_RSTIF
--   M04_CLKIF
--   M04_CLKENIF
--   S05_RSTIF
--   S05_CLKIF
--   S05_CLKENIF
--   M05_RSTIF
--   M05_CLKIF
--   M05_CLKENIF
--   S06_RSTIF
--   S06_CLKIF
--   S06_CLKENIF
--   M06_RSTIF
--   M06_CLKIF
--   M06_CLKENIF
--   S07_RSTIF
--   S07_CLKIF
--   S07_CLKENIF
--   M07_RSTIF
--   M07_CLKIF
--   M07_CLKENIF
--   S08_RSTIF
--   S08_CLKIF
--   S08_CLKENIF
--   M08_RSTIF
--   M08_CLKIF
--   M08_CLKENIF
--   S09_RSTIF
--   S09_CLKIF
--   S09_CLKENIF
--   M09_RSTIF
--   M09_CLKIF
--   M09_CLKENIF
--   S10_RSTIF
--   S10_CLKIF
--   S10_CLKENIF
--   M10_RSTIF
--   M10_CLKIF
--   M10_CLKENIF
--   S11_RSTIF
--   S11_CLKIF
--   S11_CLKENIF
--   M11_RSTIF
--   M11_CLKIF
--   M11_CLKENIF
--   S12_RSTIF
--   S12_CLKIF
--   S12_CLKENIF
--   M12_RSTIF
--   M12_CLKIF
--   M12_CLKENIF
--   S13_RSTIF
--   S13_CLKIF
--   S13_CLKENIF
--   M13_RSTIF
--   M13_CLKIF
--   M13_CLKENIF
--   S14_RSTIF
--   S14_CLKIF
--   S14_CLKENIF
--   M14_RSTIF
--   M14_CLKIF
--   M14_CLKENIF
--   S15_RSTIF
--   S15_CLKIF
--   S15_CLKENIF
--   M15_RSTIF
--   M15_CLKIF
--   M15_CLKENIF

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

LIBRARY axis_interconnect_v1_1;
USE axis_interconnect_v1_1.axis_interconnect_v1_1_axis_interconnect_16x16_top;

ENTITY axis_fifo IS
  PORT (
    ACLK : IN STD_LOGIC;
    ARESETN : IN STD_LOGIC;
    S00_AXIS_ACLK : IN STD_LOGIC;
    S00_AXIS_ARESETN : IN STD_LOGIC;
    S00_AXIS_TVALID : IN STD_LOGIC;
    S00_AXIS_TREADY : OUT STD_LOGIC;
    S00_AXIS_TDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    S00_AXIS_TLAST : IN STD_LOGIC;
    M00_AXIS_ACLK : IN STD_LOGIC;
    M00_AXIS_ARESETN : IN STD_LOGIC;
    M00_AXIS_TVALID : OUT STD_LOGIC;
    M00_AXIS_TREADY : IN STD_LOGIC;
    M00_AXIS_TDATA : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    M00_AXIS_TLAST : OUT STD_LOGIC
  );
END axis_fifo;

ARCHITECTURE spartan6 OF axis_fifo IS

  COMPONENT axis_interconnect_v1_1_axis_interconnect_16x16_top IS
    GENERIC (
      C_FAMILY : STRING;
      C_NUM_MI_SLOTS : INTEGER;
      C_NUM_SI_SLOTS : INTEGER;
      C_SWITCH_MI_REG_CONFIG : INTEGER;
      C_SWITCH_SI_REG_CONFIG : INTEGER;
      C_SWITCH_MODE : INTEGER;
      C_SWITCH_MAX_XFERS_PER_ARB : INTEGER;
      C_SWITCH_NUM_CYCLES_TIMEOUT : INTEGER;
      C_SWITCH_TDATA_WIDTH : INTEGER;
      C_SWITCH_TID_WIDTH : INTEGER;
      C_SWITCH_TDEST_WIDTH : INTEGER;
      C_SWITCH_TUSER_WIDTH : INTEGER;
      C_SWITCH_SIGNAL_SET : INTEGER;
      C_SWITCH_ACLK_RATIO : INTEGER;
      C_SWITCH_USE_ACLKEN : INTEGER;
      C_M00_AXIS_CONNECTIVITY : INTEGER;
      C_M01_AXIS_CONNECTIVITY : INTEGER;
      C_M02_AXIS_CONNECTIVITY : INTEGER;
      C_M03_AXIS_CONNECTIVITY : INTEGER;
      C_M04_AXIS_CONNECTIVITY : INTEGER;
      C_M05_AXIS_CONNECTIVITY : INTEGER;
      C_M06_AXIS_CONNECTIVITY : INTEGER;
      C_M07_AXIS_CONNECTIVITY : INTEGER;
      C_M08_AXIS_CONNECTIVITY : INTEGER;
      C_M09_AXIS_CONNECTIVITY : INTEGER;
      C_M10_AXIS_CONNECTIVITY : INTEGER;
      C_M11_AXIS_CONNECTIVITY : INTEGER;
      C_M12_AXIS_CONNECTIVITY : INTEGER;
      C_M13_AXIS_CONNECTIVITY : INTEGER;
      C_M14_AXIS_CONNECTIVITY : INTEGER;
      C_M15_AXIS_CONNECTIVITY : INTEGER;
      C_M00_AXIS_BASETDEST : INTEGER;
      C_M01_AXIS_BASETDEST : INTEGER;
      C_M02_AXIS_BASETDEST : INTEGER;
      C_M03_AXIS_BASETDEST : INTEGER;
      C_M04_AXIS_BASETDEST : INTEGER;
      C_M05_AXIS_BASETDEST : INTEGER;
      C_M06_AXIS_BASETDEST : INTEGER;
      C_M07_AXIS_BASETDEST : INTEGER;
      C_M08_AXIS_BASETDEST : INTEGER;
      C_M09_AXIS_BASETDEST : INTEGER;
      C_M10_AXIS_BASETDEST : INTEGER;
      C_M11_AXIS_BASETDEST : INTEGER;
      C_M12_AXIS_BASETDEST : INTEGER;
      C_M13_AXIS_BASETDEST : INTEGER;
      C_M14_AXIS_BASETDEST : INTEGER;
      C_M15_AXIS_BASETDEST : INTEGER;
      C_M00_AXIS_HIGHTDEST : INTEGER;
      C_M01_AXIS_HIGHTDEST : INTEGER;
      C_M02_AXIS_HIGHTDEST : INTEGER;
      C_M03_AXIS_HIGHTDEST : INTEGER;
      C_M04_AXIS_HIGHTDEST : INTEGER;
      C_M05_AXIS_HIGHTDEST : INTEGER;
      C_M06_AXIS_HIGHTDEST : INTEGER;
      C_M07_AXIS_HIGHTDEST : INTEGER;
      C_M08_AXIS_HIGHTDEST : INTEGER;
      C_M09_AXIS_HIGHTDEST : INTEGER;
      C_M10_AXIS_HIGHTDEST : INTEGER;
      C_M11_AXIS_HIGHTDEST : INTEGER;
      C_M12_AXIS_HIGHTDEST : INTEGER;
      C_M13_AXIS_HIGHTDEST : INTEGER;
      C_M14_AXIS_HIGHTDEST : INTEGER;
      C_M15_AXIS_HIGHTDEST : INTEGER;
      C_S00_AXIS_TDATA_WIDTH : INTEGER;
      C_S01_AXIS_TDATA_WIDTH : INTEGER;
      C_S02_AXIS_TDATA_WIDTH : INTEGER;
      C_S03_AXIS_TDATA_WIDTH : INTEGER;
      C_S04_AXIS_TDATA_WIDTH : INTEGER;
      C_S05_AXIS_TDATA_WIDTH : INTEGER;
      C_S06_AXIS_TDATA_WIDTH : INTEGER;
      C_S07_AXIS_TDATA_WIDTH : INTEGER;
      C_S08_AXIS_TDATA_WIDTH : INTEGER;
      C_S09_AXIS_TDATA_WIDTH : INTEGER;
      C_S10_AXIS_TDATA_WIDTH : INTEGER;
      C_S11_AXIS_TDATA_WIDTH : INTEGER;
      C_S12_AXIS_TDATA_WIDTH : INTEGER;
      C_S13_AXIS_TDATA_WIDTH : INTEGER;
      C_S14_AXIS_TDATA_WIDTH : INTEGER;
      C_S15_AXIS_TDATA_WIDTH : INTEGER;
      C_S00_AXIS_TUSER_WIDTH : INTEGER;
      C_S01_AXIS_TUSER_WIDTH : INTEGER;
      C_S02_AXIS_TUSER_WIDTH : INTEGER;
      C_S03_AXIS_TUSER_WIDTH : INTEGER;
      C_S04_AXIS_TUSER_WIDTH : INTEGER;
      C_S05_AXIS_TUSER_WIDTH : INTEGER;
      C_S06_AXIS_TUSER_WIDTH : INTEGER;
      C_S07_AXIS_TUSER_WIDTH : INTEGER;
      C_S08_AXIS_TUSER_WIDTH : INTEGER;
      C_S09_AXIS_TUSER_WIDTH : INTEGER;
      C_S10_AXIS_TUSER_WIDTH : INTEGER;
      C_S11_AXIS_TUSER_WIDTH : INTEGER;
      C_S12_AXIS_TUSER_WIDTH : INTEGER;
      C_S13_AXIS_TUSER_WIDTH : INTEGER;
      C_S14_AXIS_TUSER_WIDTH : INTEGER;
      C_S15_AXIS_TUSER_WIDTH : INTEGER;
      C_S00_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_S01_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_S02_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_S03_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_S04_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_S05_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_S06_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_S07_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_S08_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_S09_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_S10_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_S11_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_S12_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_S13_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_S14_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_S15_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_S00_AXIS_ACLK_RATIO : INTEGER;
      C_S01_AXIS_ACLK_RATIO : INTEGER;
      C_S02_AXIS_ACLK_RATIO : INTEGER;
      C_S03_AXIS_ACLK_RATIO : INTEGER;
      C_S04_AXIS_ACLK_RATIO : INTEGER;
      C_S05_AXIS_ACLK_RATIO : INTEGER;
      C_S06_AXIS_ACLK_RATIO : INTEGER;
      C_S07_AXIS_ACLK_RATIO : INTEGER;
      C_S08_AXIS_ACLK_RATIO : INTEGER;
      C_S09_AXIS_ACLK_RATIO : INTEGER;
      C_S10_AXIS_ACLK_RATIO : INTEGER;
      C_S11_AXIS_ACLK_RATIO : INTEGER;
      C_S12_AXIS_ACLK_RATIO : INTEGER;
      C_S13_AXIS_ACLK_RATIO : INTEGER;
      C_S14_AXIS_ACLK_RATIO : INTEGER;
      C_S15_AXIS_ACLK_RATIO : INTEGER;
      C_S00_AXIS_REG_CONFIG : INTEGER;
      C_S01_AXIS_REG_CONFIG : INTEGER;
      C_S02_AXIS_REG_CONFIG : INTEGER;
      C_S03_AXIS_REG_CONFIG : INTEGER;
      C_S04_AXIS_REG_CONFIG : INTEGER;
      C_S05_AXIS_REG_CONFIG : INTEGER;
      C_S06_AXIS_REG_CONFIG : INTEGER;
      C_S07_AXIS_REG_CONFIG : INTEGER;
      C_S08_AXIS_REG_CONFIG : INTEGER;
      C_S09_AXIS_REG_CONFIG : INTEGER;
      C_S10_AXIS_REG_CONFIG : INTEGER;
      C_S11_AXIS_REG_CONFIG : INTEGER;
      C_S12_AXIS_REG_CONFIG : INTEGER;
      C_S13_AXIS_REG_CONFIG : INTEGER;
      C_S14_AXIS_REG_CONFIG : INTEGER;
      C_S15_AXIS_REG_CONFIG : INTEGER;
      C_S00_AXIS_FIFO_DEPTH : INTEGER;
      C_S01_AXIS_FIFO_DEPTH : INTEGER;
      C_S02_AXIS_FIFO_DEPTH : INTEGER;
      C_S03_AXIS_FIFO_DEPTH : INTEGER;
      C_S04_AXIS_FIFO_DEPTH : INTEGER;
      C_S05_AXIS_FIFO_DEPTH : INTEGER;
      C_S06_AXIS_FIFO_DEPTH : INTEGER;
      C_S07_AXIS_FIFO_DEPTH : INTEGER;
      C_S08_AXIS_FIFO_DEPTH : INTEGER;
      C_S09_AXIS_FIFO_DEPTH : INTEGER;
      C_S10_AXIS_FIFO_DEPTH : INTEGER;
      C_S11_AXIS_FIFO_DEPTH : INTEGER;
      C_S12_AXIS_FIFO_DEPTH : INTEGER;
      C_S13_AXIS_FIFO_DEPTH : INTEGER;
      C_S14_AXIS_FIFO_DEPTH : INTEGER;
      C_S15_AXIS_FIFO_DEPTH : INTEGER;
      C_S00_AXIS_FIFO_MODE : INTEGER;
      C_S01_AXIS_FIFO_MODE : INTEGER;
      C_S02_AXIS_FIFO_MODE : INTEGER;
      C_S03_AXIS_FIFO_MODE : INTEGER;
      C_S04_AXIS_FIFO_MODE : INTEGER;
      C_S05_AXIS_FIFO_MODE : INTEGER;
      C_S06_AXIS_FIFO_MODE : INTEGER;
      C_S07_AXIS_FIFO_MODE : INTEGER;
      C_S08_AXIS_FIFO_MODE : INTEGER;
      C_S09_AXIS_FIFO_MODE : INTEGER;
      C_S10_AXIS_FIFO_MODE : INTEGER;
      C_S11_AXIS_FIFO_MODE : INTEGER;
      C_S12_AXIS_FIFO_MODE : INTEGER;
      C_S13_AXIS_FIFO_MODE : INTEGER;
      C_S14_AXIS_FIFO_MODE : INTEGER;
      C_S15_AXIS_FIFO_MODE : INTEGER;
      C_M00_AXIS_TDATA_WIDTH : INTEGER;
      C_M01_AXIS_TDATA_WIDTH : INTEGER;
      C_M02_AXIS_TDATA_WIDTH : INTEGER;
      C_M03_AXIS_TDATA_WIDTH : INTEGER;
      C_M04_AXIS_TDATA_WIDTH : INTEGER;
      C_M05_AXIS_TDATA_WIDTH : INTEGER;
      C_M06_AXIS_TDATA_WIDTH : INTEGER;
      C_M07_AXIS_TDATA_WIDTH : INTEGER;
      C_M08_AXIS_TDATA_WIDTH : INTEGER;
      C_M09_AXIS_TDATA_WIDTH : INTEGER;
      C_M10_AXIS_TDATA_WIDTH : INTEGER;
      C_M11_AXIS_TDATA_WIDTH : INTEGER;
      C_M12_AXIS_TDATA_WIDTH : INTEGER;
      C_M13_AXIS_TDATA_WIDTH : INTEGER;
      C_M14_AXIS_TDATA_WIDTH : INTEGER;
      C_M15_AXIS_TDATA_WIDTH : INTEGER;
      C_M00_AXIS_TUSER_WIDTH : INTEGER;
      C_M01_AXIS_TUSER_WIDTH : INTEGER;
      C_M02_AXIS_TUSER_WIDTH : INTEGER;
      C_M03_AXIS_TUSER_WIDTH : INTEGER;
      C_M04_AXIS_TUSER_WIDTH : INTEGER;
      C_M05_AXIS_TUSER_WIDTH : INTEGER;
      C_M06_AXIS_TUSER_WIDTH : INTEGER;
      C_M07_AXIS_TUSER_WIDTH : INTEGER;
      C_M08_AXIS_TUSER_WIDTH : INTEGER;
      C_M09_AXIS_TUSER_WIDTH : INTEGER;
      C_M10_AXIS_TUSER_WIDTH : INTEGER;
      C_M11_AXIS_TUSER_WIDTH : INTEGER;
      C_M12_AXIS_TUSER_WIDTH : INTEGER;
      C_M13_AXIS_TUSER_WIDTH : INTEGER;
      C_M14_AXIS_TUSER_WIDTH : INTEGER;
      C_M15_AXIS_TUSER_WIDTH : INTEGER;
      C_M00_AXIS_ACLK_RATIO : INTEGER;
      C_M01_AXIS_ACLK_RATIO : INTEGER;
      C_M02_AXIS_ACLK_RATIO : INTEGER;
      C_M03_AXIS_ACLK_RATIO : INTEGER;
      C_M04_AXIS_ACLK_RATIO : INTEGER;
      C_M05_AXIS_ACLK_RATIO : INTEGER;
      C_M06_AXIS_ACLK_RATIO : INTEGER;
      C_M07_AXIS_ACLK_RATIO : INTEGER;
      C_M08_AXIS_ACLK_RATIO : INTEGER;
      C_M09_AXIS_ACLK_RATIO : INTEGER;
      C_M10_AXIS_ACLK_RATIO : INTEGER;
      C_M11_AXIS_ACLK_RATIO : INTEGER;
      C_M12_AXIS_ACLK_RATIO : INTEGER;
      C_M13_AXIS_ACLK_RATIO : INTEGER;
      C_M14_AXIS_ACLK_RATIO : INTEGER;
      C_M15_AXIS_ACLK_RATIO : INTEGER;
      C_M00_AXIS_REG_CONFIG : INTEGER;
      C_M01_AXIS_REG_CONFIG : INTEGER;
      C_M02_AXIS_REG_CONFIG : INTEGER;
      C_M03_AXIS_REG_CONFIG : INTEGER;
      C_M04_AXIS_REG_CONFIG : INTEGER;
      C_M05_AXIS_REG_CONFIG : INTEGER;
      C_M06_AXIS_REG_CONFIG : INTEGER;
      C_M07_AXIS_REG_CONFIG : INTEGER;
      C_M08_AXIS_REG_CONFIG : INTEGER;
      C_M09_AXIS_REG_CONFIG : INTEGER;
      C_M10_AXIS_REG_CONFIG : INTEGER;
      C_M11_AXIS_REG_CONFIG : INTEGER;
      C_M12_AXIS_REG_CONFIG : INTEGER;
      C_M13_AXIS_REG_CONFIG : INTEGER;
      C_M14_AXIS_REG_CONFIG : INTEGER;
      C_M15_AXIS_REG_CONFIG : INTEGER;
      C_M00_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_M01_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_M02_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_M03_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_M04_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_M05_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_M06_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_M07_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_M08_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_M09_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_M10_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_M11_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_M12_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_M13_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_M14_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_M15_AXIS_IS_ACLK_ASYNC : INTEGER;
      C_M00_AXIS_FIFO_DEPTH : INTEGER;
      C_M01_AXIS_FIFO_DEPTH : INTEGER;
      C_M02_AXIS_FIFO_DEPTH : INTEGER;
      C_M03_AXIS_FIFO_DEPTH : INTEGER;
      C_M04_AXIS_FIFO_DEPTH : INTEGER;
      C_M05_AXIS_FIFO_DEPTH : INTEGER;
      C_M06_AXIS_FIFO_DEPTH : INTEGER;
      C_M07_AXIS_FIFO_DEPTH : INTEGER;
      C_M08_AXIS_FIFO_DEPTH : INTEGER;
      C_M09_AXIS_FIFO_DEPTH : INTEGER;
      C_M10_AXIS_FIFO_DEPTH : INTEGER;
      C_M11_AXIS_FIFO_DEPTH : INTEGER;
      C_M12_AXIS_FIFO_DEPTH : INTEGER;
      C_M13_AXIS_FIFO_DEPTH : INTEGER;
      C_M14_AXIS_FIFO_DEPTH : INTEGER;
      C_M15_AXIS_FIFO_DEPTH : INTEGER;
      C_M00_AXIS_FIFO_MODE : INTEGER;
      C_M01_AXIS_FIFO_MODE : INTEGER;
      C_M02_AXIS_FIFO_MODE : INTEGER;
      C_M03_AXIS_FIFO_MODE : INTEGER;
      C_M04_AXIS_FIFO_MODE : INTEGER;
      C_M05_AXIS_FIFO_MODE : INTEGER;
      C_M06_AXIS_FIFO_MODE : INTEGER;
      C_M07_AXIS_FIFO_MODE : INTEGER;
      C_M08_AXIS_FIFO_MODE : INTEGER;
      C_M09_AXIS_FIFO_MODE : INTEGER;
      C_M10_AXIS_FIFO_MODE : INTEGER;
      C_M11_AXIS_FIFO_MODE : INTEGER;
      C_M12_AXIS_FIFO_MODE : INTEGER;
      C_M13_AXIS_FIFO_MODE : INTEGER;
      C_M14_AXIS_FIFO_MODE : INTEGER;
      C_M15_AXIS_FIFO_MODE : INTEGER
    );
    PORT (
      ACLK : IN STD_LOGIC;
      ARESETN : IN STD_LOGIC;
      S00_AXIS_ACLK : IN STD_LOGIC;
      S00_AXIS_ARESETN : IN STD_LOGIC;
      S00_AXIS_TVALID : IN STD_LOGIC;
      S00_AXIS_TREADY : OUT STD_LOGIC;
      S00_AXIS_TDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      S00_AXIS_TLAST : IN STD_LOGIC;
      M00_AXIS_ACLK : IN STD_LOGIC;
      M00_AXIS_ARESETN : IN STD_LOGIC;
      M00_AXIS_TVALID : OUT STD_LOGIC;
      M00_AXIS_TREADY : IN STD_LOGIC;
      M00_AXIS_TDATA : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
      M00_AXIS_TLAST : OUT STD_LOGIC;
      ACLKEN : IN STD_LOGIC;
      S01_AXIS_ACLK : IN STD_LOGIC;
      S02_AXIS_ACLK : IN STD_LOGIC;
      S03_AXIS_ACLK : IN STD_LOGIC;
      S04_AXIS_ACLK : IN STD_LOGIC;
      S05_AXIS_ACLK : IN STD_LOGIC;
      S06_AXIS_ACLK : IN STD_LOGIC;
      S07_AXIS_ACLK : IN STD_LOGIC;
      S08_AXIS_ACLK : IN STD_LOGIC;
      S09_AXIS_ACLK : IN STD_LOGIC;
      S10_AXIS_ACLK : IN STD_LOGIC;
      S11_AXIS_ACLK : IN STD_LOGIC;
      S12_AXIS_ACLK : IN STD_LOGIC;
      S13_AXIS_ACLK : IN STD_LOGIC;
      S14_AXIS_ACLK : IN STD_LOGIC;
      S15_AXIS_ACLK : IN STD_LOGIC;
      S01_AXIS_ARESETN : IN STD_LOGIC;
      S02_AXIS_ARESETN : IN STD_LOGIC;
      S03_AXIS_ARESETN : IN STD_LOGIC;
      S04_AXIS_ARESETN : IN STD_LOGIC;
      S05_AXIS_ARESETN : IN STD_LOGIC;
      S06_AXIS_ARESETN : IN STD_LOGIC;
      S07_AXIS_ARESETN : IN STD_LOGIC;
      S08_AXIS_ARESETN : IN STD_LOGIC;
      S09_AXIS_ARESETN : IN STD_LOGIC;
      S10_AXIS_ARESETN : IN STD_LOGIC;
      S11_AXIS_ARESETN : IN STD_LOGIC;
      S12_AXIS_ARESETN : IN STD_LOGIC;
      S13_AXIS_ARESETN : IN STD_LOGIC;
      S14_AXIS_ARESETN : IN STD_LOGIC;
      S15_AXIS_ARESETN : IN STD_LOGIC;
      S00_AXIS_ACLKEN : IN STD_LOGIC;
      S01_AXIS_ACLKEN : IN STD_LOGIC;
      S02_AXIS_ACLKEN : IN STD_LOGIC;
      S03_AXIS_ACLKEN : IN STD_LOGIC;
      S04_AXIS_ACLKEN : IN STD_LOGIC;
      S05_AXIS_ACLKEN : IN STD_LOGIC;
      S06_AXIS_ACLKEN : IN STD_LOGIC;
      S07_AXIS_ACLKEN : IN STD_LOGIC;
      S08_AXIS_ACLKEN : IN STD_LOGIC;
      S09_AXIS_ACLKEN : IN STD_LOGIC;
      S10_AXIS_ACLKEN : IN STD_LOGIC;
      S11_AXIS_ACLKEN : IN STD_LOGIC;
      S12_AXIS_ACLKEN : IN STD_LOGIC;
      S13_AXIS_ACLKEN : IN STD_LOGIC;
      S14_AXIS_ACLKEN : IN STD_LOGIC;
      S15_AXIS_ACLKEN : IN STD_LOGIC;
      S01_AXIS_TVALID : IN STD_LOGIC;
      S02_AXIS_TVALID : IN STD_LOGIC;
      S03_AXIS_TVALID : IN STD_LOGIC;
      S04_AXIS_TVALID : IN STD_LOGIC;
      S05_AXIS_TVALID : IN STD_LOGIC;
      S06_AXIS_TVALID : IN STD_LOGIC;
      S07_AXIS_TVALID : IN STD_LOGIC;
      S08_AXIS_TVALID : IN STD_LOGIC;
      S09_AXIS_TVALID : IN STD_LOGIC;
      S10_AXIS_TVALID : IN STD_LOGIC;
      S11_AXIS_TVALID : IN STD_LOGIC;
      S12_AXIS_TVALID : IN STD_LOGIC;
      S13_AXIS_TVALID : IN STD_LOGIC;
      S14_AXIS_TVALID : IN STD_LOGIC;
      S15_AXIS_TVALID : IN STD_LOGIC;
      S01_AXIS_TDATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S02_AXIS_TDATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S03_AXIS_TDATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S04_AXIS_TDATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S05_AXIS_TDATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S06_AXIS_TDATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S07_AXIS_TDATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S08_AXIS_TDATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S09_AXIS_TDATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S10_AXIS_TDATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S11_AXIS_TDATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S12_AXIS_TDATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S13_AXIS_TDATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S14_AXIS_TDATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S15_AXIS_TDATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      S00_AXIS_TSTRB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S01_AXIS_TSTRB : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S02_AXIS_TSTRB : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S03_AXIS_TSTRB : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S04_AXIS_TSTRB : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S05_AXIS_TSTRB : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S06_AXIS_TSTRB : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S07_AXIS_TSTRB : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S08_AXIS_TSTRB : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S09_AXIS_TSTRB : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S10_AXIS_TSTRB : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S11_AXIS_TSTRB : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S12_AXIS_TSTRB : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S13_AXIS_TSTRB : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S14_AXIS_TSTRB : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S15_AXIS_TSTRB : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S00_AXIS_TKEEP : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S01_AXIS_TKEEP : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S02_AXIS_TKEEP : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S03_AXIS_TKEEP : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S04_AXIS_TKEEP : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S05_AXIS_TKEEP : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S06_AXIS_TKEEP : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S07_AXIS_TKEEP : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S08_AXIS_TKEEP : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S09_AXIS_TKEEP : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S10_AXIS_TKEEP : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S11_AXIS_TKEEP : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S12_AXIS_TKEEP : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S13_AXIS_TKEEP : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S14_AXIS_TKEEP : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S15_AXIS_TKEEP : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S01_AXIS_TLAST : IN STD_LOGIC;
      S02_AXIS_TLAST : IN STD_LOGIC;
      S03_AXIS_TLAST : IN STD_LOGIC;
      S04_AXIS_TLAST : IN STD_LOGIC;
      S05_AXIS_TLAST : IN STD_LOGIC;
      S06_AXIS_TLAST : IN STD_LOGIC;
      S07_AXIS_TLAST : IN STD_LOGIC;
      S08_AXIS_TLAST : IN STD_LOGIC;
      S09_AXIS_TLAST : IN STD_LOGIC;
      S10_AXIS_TLAST : IN STD_LOGIC;
      S11_AXIS_TLAST : IN STD_LOGIC;
      S12_AXIS_TLAST : IN STD_LOGIC;
      S13_AXIS_TLAST : IN STD_LOGIC;
      S14_AXIS_TLAST : IN STD_LOGIC;
      S15_AXIS_TLAST : IN STD_LOGIC;
      S00_AXIS_TID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S01_AXIS_TID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S02_AXIS_TID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S03_AXIS_TID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S04_AXIS_TID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S05_AXIS_TID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S06_AXIS_TID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S07_AXIS_TID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S08_AXIS_TID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S09_AXIS_TID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S10_AXIS_TID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S11_AXIS_TID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S12_AXIS_TID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S13_AXIS_TID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S14_AXIS_TID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S15_AXIS_TID : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S00_AXIS_TDEST : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S01_AXIS_TDEST : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S02_AXIS_TDEST : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S03_AXIS_TDEST : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S04_AXIS_TDEST : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S05_AXIS_TDEST : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S06_AXIS_TDEST : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S07_AXIS_TDEST : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S08_AXIS_TDEST : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S09_AXIS_TDEST : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S10_AXIS_TDEST : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S11_AXIS_TDEST : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S12_AXIS_TDEST : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S13_AXIS_TDEST : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S14_AXIS_TDEST : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S15_AXIS_TDEST : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S00_AXIS_TUSER : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      S01_AXIS_TUSER : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S02_AXIS_TUSER : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S03_AXIS_TUSER : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S04_AXIS_TUSER : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S05_AXIS_TUSER : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S06_AXIS_TUSER : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S07_AXIS_TUSER : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S08_AXIS_TUSER : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S09_AXIS_TUSER : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S10_AXIS_TUSER : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S11_AXIS_TUSER : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S12_AXIS_TUSER : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S13_AXIS_TUSER : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S14_AXIS_TUSER : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      S15_AXIS_TUSER : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      M01_AXIS_ACLK : IN STD_LOGIC;
      M02_AXIS_ACLK : IN STD_LOGIC;
      M03_AXIS_ACLK : IN STD_LOGIC;
      M04_AXIS_ACLK : IN STD_LOGIC;
      M05_AXIS_ACLK : IN STD_LOGIC;
      M06_AXIS_ACLK : IN STD_LOGIC;
      M07_AXIS_ACLK : IN STD_LOGIC;
      M08_AXIS_ACLK : IN STD_LOGIC;
      M09_AXIS_ACLK : IN STD_LOGIC;
      M10_AXIS_ACLK : IN STD_LOGIC;
      M11_AXIS_ACLK : IN STD_LOGIC;
      M12_AXIS_ACLK : IN STD_LOGIC;
      M13_AXIS_ACLK : IN STD_LOGIC;
      M14_AXIS_ACLK : IN STD_LOGIC;
      M15_AXIS_ACLK : IN STD_LOGIC;
      M01_AXIS_ARESETN : IN STD_LOGIC;
      M02_AXIS_ARESETN : IN STD_LOGIC;
      M03_AXIS_ARESETN : IN STD_LOGIC;
      M04_AXIS_ARESETN : IN STD_LOGIC;
      M05_AXIS_ARESETN : IN STD_LOGIC;
      M06_AXIS_ARESETN : IN STD_LOGIC;
      M07_AXIS_ARESETN : IN STD_LOGIC;
      M08_AXIS_ARESETN : IN STD_LOGIC;
      M09_AXIS_ARESETN : IN STD_LOGIC;
      M10_AXIS_ARESETN : IN STD_LOGIC;
      M11_AXIS_ARESETN : IN STD_LOGIC;
      M12_AXIS_ARESETN : IN STD_LOGIC;
      M13_AXIS_ARESETN : IN STD_LOGIC;
      M14_AXIS_ARESETN : IN STD_LOGIC;
      M15_AXIS_ARESETN : IN STD_LOGIC;
      M00_AXIS_ACLKEN : IN STD_LOGIC;
      M01_AXIS_ACLKEN : IN STD_LOGIC;
      M02_AXIS_ACLKEN : IN STD_LOGIC;
      M03_AXIS_ACLKEN : IN STD_LOGIC;
      M04_AXIS_ACLKEN : IN STD_LOGIC;
      M05_AXIS_ACLKEN : IN STD_LOGIC;
      M06_AXIS_ACLKEN : IN STD_LOGIC;
      M07_AXIS_ACLKEN : IN STD_LOGIC;
      M08_AXIS_ACLKEN : IN STD_LOGIC;
      M09_AXIS_ACLKEN : IN STD_LOGIC;
      M10_AXIS_ACLKEN : IN STD_LOGIC;
      M11_AXIS_ACLKEN : IN STD_LOGIC;
      M12_AXIS_ACLKEN : IN STD_LOGIC;
      M13_AXIS_ACLKEN : IN STD_LOGIC;
      M14_AXIS_ACLKEN : IN STD_LOGIC;
      M15_AXIS_ACLKEN : IN STD_LOGIC;
      M01_AXIS_TREADY : IN STD_LOGIC;
      M02_AXIS_TREADY : IN STD_LOGIC;
      M03_AXIS_TREADY : IN STD_LOGIC;
      M04_AXIS_TREADY : IN STD_LOGIC;
      M05_AXIS_TREADY : IN STD_LOGIC;
      M06_AXIS_TREADY : IN STD_LOGIC;
      M07_AXIS_TREADY : IN STD_LOGIC;
      M08_AXIS_TREADY : IN STD_LOGIC;
      M09_AXIS_TREADY : IN STD_LOGIC;
      M10_AXIS_TREADY : IN STD_LOGIC;
      M11_AXIS_TREADY : IN STD_LOGIC;
      M12_AXIS_TREADY : IN STD_LOGIC;
      M13_AXIS_TREADY : IN STD_LOGIC;
      M14_AXIS_TREADY : IN STD_LOGIC;
      M15_AXIS_TREADY : IN STD_LOGIC;
      S00_ARB_REQ_SUPPRESS : IN STD_LOGIC;
      S01_ARB_REQ_SUPPRESS : IN STD_LOGIC;
      S02_ARB_REQ_SUPPRESS : IN STD_LOGIC;
      S03_ARB_REQ_SUPPRESS : IN STD_LOGIC;
      S04_ARB_REQ_SUPPRESS : IN STD_LOGIC;
      S05_ARB_REQ_SUPPRESS : IN STD_LOGIC;
      S06_ARB_REQ_SUPPRESS : IN STD_LOGIC;
      S07_ARB_REQ_SUPPRESS : IN STD_LOGIC;
      S08_ARB_REQ_SUPPRESS : IN STD_LOGIC;
      S09_ARB_REQ_SUPPRESS : IN STD_LOGIC;
      S10_ARB_REQ_SUPPRESS : IN STD_LOGIC;
      S11_ARB_REQ_SUPPRESS : IN STD_LOGIC;
      S12_ARB_REQ_SUPPRESS : IN STD_LOGIC;
      S13_ARB_REQ_SUPPRESS : IN STD_LOGIC;
      S14_ARB_REQ_SUPPRESS : IN STD_LOGIC;
      S15_ARB_REQ_SUPPRESS : IN STD_LOGIC
    );
  END COMPONENT axis_interconnect_v1_1_axis_interconnect_16x16_top;

BEGIN

  U0 : axis_interconnect_v1_1_axis_interconnect_16x16_top
    GENERIC MAP (
      C_FAMILY => "spartan6",
      C_M00_AXIS_ACLK_RATIO => 12,
      C_M00_AXIS_BASETDEST => X"0",
      C_M00_AXIS_CONNECTIVITY => X"FFFF",
      C_M00_AXIS_FIFO_DEPTH => 32,
      C_M00_AXIS_FIFO_MODE => 0,
      C_M00_AXIS_HIGHTDEST => X"0",
      C_M00_AXIS_IS_ACLK_ASYNC => 0,
      C_M00_AXIS_REG_CONFIG => 0,
      C_M00_AXIS_TDATA_WIDTH => 8,
      C_M00_AXIS_TUSER_WIDTH => 1,
      C_M01_AXIS_ACLK_RATIO => 12,
      C_M01_AXIS_BASETDEST => X"1",
      C_M01_AXIS_CONNECTIVITY => X"FFFF",
      C_M01_AXIS_FIFO_DEPTH => 32,
      C_M01_AXIS_FIFO_MODE => 0,
      C_M01_AXIS_HIGHTDEST => X"1",
      C_M01_AXIS_IS_ACLK_ASYNC => 0,
      C_M01_AXIS_REG_CONFIG => 0,
      C_M01_AXIS_TDATA_WIDTH => 8,
      C_M01_AXIS_TUSER_WIDTH => 1,
      C_M02_AXIS_ACLK_RATIO => 12,
      C_M02_AXIS_BASETDEST => X"2",
      C_M02_AXIS_CONNECTIVITY => X"FFFF",
      C_M02_AXIS_FIFO_DEPTH => 32,
      C_M02_AXIS_FIFO_MODE => 0,
      C_M02_AXIS_HIGHTDEST => X"2",
      C_M02_AXIS_IS_ACLK_ASYNC => 0,
      C_M02_AXIS_REG_CONFIG => 0,
      C_M02_AXIS_TDATA_WIDTH => 8,
      C_M02_AXIS_TUSER_WIDTH => 1,
      C_M03_AXIS_ACLK_RATIO => 12,
      C_M03_AXIS_BASETDEST => X"3",
      C_M03_AXIS_CONNECTIVITY => X"FFFF",
      C_M03_AXIS_FIFO_DEPTH => 32,
      C_M03_AXIS_FIFO_MODE => 0,
      C_M03_AXIS_HIGHTDEST => X"3",
      C_M03_AXIS_IS_ACLK_ASYNC => 0,
      C_M03_AXIS_REG_CONFIG => 0,
      C_M03_AXIS_TDATA_WIDTH => 8,
      C_M03_AXIS_TUSER_WIDTH => 1,
      C_M04_AXIS_ACLK_RATIO => 12,
      C_M04_AXIS_BASETDEST => X"4",
      C_M04_AXIS_CONNECTIVITY => X"FFFF",
      C_M04_AXIS_FIFO_DEPTH => 32,
      C_M04_AXIS_FIFO_MODE => 0,
      C_M04_AXIS_HIGHTDEST => X"4",
      C_M04_AXIS_IS_ACLK_ASYNC => 0,
      C_M04_AXIS_REG_CONFIG => 0,
      C_M04_AXIS_TDATA_WIDTH => 8,
      C_M04_AXIS_TUSER_WIDTH => 1,
      C_M05_AXIS_ACLK_RATIO => 12,
      C_M05_AXIS_BASETDEST => X"5",
      C_M05_AXIS_CONNECTIVITY => X"FFFF",
      C_M05_AXIS_FIFO_DEPTH => 32,
      C_M05_AXIS_FIFO_MODE => 0,
      C_M05_AXIS_HIGHTDEST => X"5",
      C_M05_AXIS_IS_ACLK_ASYNC => 0,
      C_M05_AXIS_REG_CONFIG => 0,
      C_M05_AXIS_TDATA_WIDTH => 8,
      C_M05_AXIS_TUSER_WIDTH => 1,
      C_M06_AXIS_ACLK_RATIO => 12,
      C_M06_AXIS_BASETDEST => X"6",
      C_M06_AXIS_CONNECTIVITY => X"FFFF",
      C_M06_AXIS_FIFO_DEPTH => 32,
      C_M06_AXIS_FIFO_MODE => 0,
      C_M06_AXIS_HIGHTDEST => X"6",
      C_M06_AXIS_IS_ACLK_ASYNC => 0,
      C_M06_AXIS_REG_CONFIG => 0,
      C_M06_AXIS_TDATA_WIDTH => 8,
      C_M06_AXIS_TUSER_WIDTH => 1,
      C_M07_AXIS_ACLK_RATIO => 12,
      C_M07_AXIS_BASETDEST => X"7",
      C_M07_AXIS_CONNECTIVITY => X"FFFF",
      C_M07_AXIS_FIFO_DEPTH => 32,
      C_M07_AXIS_FIFO_MODE => 0,
      C_M07_AXIS_HIGHTDEST => X"7",
      C_M07_AXIS_IS_ACLK_ASYNC => 0,
      C_M07_AXIS_REG_CONFIG => 0,
      C_M07_AXIS_TDATA_WIDTH => 8,
      C_M07_AXIS_TUSER_WIDTH => 1,
      C_M08_AXIS_ACLK_RATIO => 12,
      C_M08_AXIS_BASETDEST => X"8",
      C_M08_AXIS_CONNECTIVITY => X"FFFF",
      C_M08_AXIS_FIFO_DEPTH => 32,
      C_M08_AXIS_FIFO_MODE => 0,
      C_M08_AXIS_HIGHTDEST => X"8",
      C_M08_AXIS_IS_ACLK_ASYNC => 0,
      C_M08_AXIS_REG_CONFIG => 0,
      C_M08_AXIS_TDATA_WIDTH => 8,
      C_M08_AXIS_TUSER_WIDTH => 1,
      C_M09_AXIS_ACLK_RATIO => 12,
      C_M09_AXIS_BASETDEST => X"9",
      C_M09_AXIS_CONNECTIVITY => X"FFFF",
      C_M09_AXIS_FIFO_DEPTH => 32,
      C_M09_AXIS_FIFO_MODE => 0,
      C_M09_AXIS_HIGHTDEST => X"9",
      C_M09_AXIS_IS_ACLK_ASYNC => 0,
      C_M09_AXIS_REG_CONFIG => 0,
      C_M09_AXIS_TDATA_WIDTH => 8,
      C_M09_AXIS_TUSER_WIDTH => 1,
      C_M10_AXIS_ACLK_RATIO => 12,
      C_M10_AXIS_BASETDEST => X"A",
      C_M10_AXIS_CONNECTIVITY => X"FFFF",
      C_M10_AXIS_FIFO_DEPTH => 32,
      C_M10_AXIS_FIFO_MODE => 0,
      C_M10_AXIS_HIGHTDEST => X"A",
      C_M10_AXIS_IS_ACLK_ASYNC => 0,
      C_M10_AXIS_REG_CONFIG => 0,
      C_M10_AXIS_TDATA_WIDTH => 8,
      C_M10_AXIS_TUSER_WIDTH => 1,
      C_M11_AXIS_ACLK_RATIO => 12,
      C_M11_AXIS_BASETDEST => X"B",
      C_M11_AXIS_CONNECTIVITY => X"FFFF",
      C_M11_AXIS_FIFO_DEPTH => 32,
      C_M11_AXIS_FIFO_MODE => 0,
      C_M11_AXIS_HIGHTDEST => X"B",
      C_M11_AXIS_IS_ACLK_ASYNC => 0,
      C_M11_AXIS_REG_CONFIG => 0,
      C_M11_AXIS_TDATA_WIDTH => 8,
      C_M11_AXIS_TUSER_WIDTH => 1,
      C_M12_AXIS_ACLK_RATIO => 12,
      C_M12_AXIS_BASETDEST => X"C",
      C_M12_AXIS_CONNECTIVITY => X"FFFF",
      C_M12_AXIS_FIFO_DEPTH => 32,
      C_M12_AXIS_FIFO_MODE => 0,
      C_M12_AXIS_HIGHTDEST => X"C",
      C_M12_AXIS_IS_ACLK_ASYNC => 0,
      C_M12_AXIS_REG_CONFIG => 0,
      C_M12_AXIS_TDATA_WIDTH => 8,
      C_M12_AXIS_TUSER_WIDTH => 1,
      C_M13_AXIS_ACLK_RATIO => 12,
      C_M13_AXIS_BASETDEST => X"D",
      C_M13_AXIS_CONNECTIVITY => X"FFFF",
      C_M13_AXIS_FIFO_DEPTH => 32,
      C_M13_AXIS_FIFO_MODE => 0,
      C_M13_AXIS_HIGHTDEST => X"D",
      C_M13_AXIS_IS_ACLK_ASYNC => 0,
      C_M13_AXIS_REG_CONFIG => 0,
      C_M13_AXIS_TDATA_WIDTH => 8,
      C_M13_AXIS_TUSER_WIDTH => 1,
      C_M14_AXIS_ACLK_RATIO => 12,
      C_M14_AXIS_BASETDEST => X"E",
      C_M14_AXIS_CONNECTIVITY => X"FFFF",
      C_M14_AXIS_FIFO_DEPTH => 32,
      C_M14_AXIS_FIFO_MODE => 0,
      C_M14_AXIS_HIGHTDEST => X"E",
      C_M14_AXIS_IS_ACLK_ASYNC => 0,
      C_M14_AXIS_REG_CONFIG => 0,
      C_M14_AXIS_TDATA_WIDTH => 8,
      C_M14_AXIS_TUSER_WIDTH => 1,
      C_M15_AXIS_ACLK_RATIO => 12,
      C_M15_AXIS_BASETDEST => X"F",
      C_M15_AXIS_CONNECTIVITY => X"FFFF",
      C_M15_AXIS_FIFO_DEPTH => 32,
      C_M15_AXIS_FIFO_MODE => 0,
      C_M15_AXIS_HIGHTDEST => X"F",
      C_M15_AXIS_IS_ACLK_ASYNC => 0,
      C_M15_AXIS_REG_CONFIG => 0,
      C_M15_AXIS_TDATA_WIDTH => 8,
      C_M15_AXIS_TUSER_WIDTH => 1,
      C_NUM_MI_SLOTS => 1,
      C_NUM_SI_SLOTS => 1,
      C_S00_AXIS_ACLK_RATIO => 12,
      C_S00_AXIS_FIFO_DEPTH => 32,
      C_S00_AXIS_FIFO_MODE => 0,
      C_S00_AXIS_IS_ACLK_ASYNC => 0,
      C_S00_AXIS_REG_CONFIG => 0,
      C_S00_AXIS_TDATA_WIDTH => 32,
      C_S00_AXIS_TUSER_WIDTH => 4,
      C_S01_AXIS_ACLK_RATIO => 12,
      C_S01_AXIS_FIFO_DEPTH => 32,
      C_S01_AXIS_FIFO_MODE => 0,
      C_S01_AXIS_IS_ACLK_ASYNC => 0,
      C_S01_AXIS_REG_CONFIG => 0,
      C_S01_AXIS_TDATA_WIDTH => 8,
      C_S01_AXIS_TUSER_WIDTH => 1,
      C_S02_AXIS_ACLK_RATIO => 12,
      C_S02_AXIS_FIFO_DEPTH => 32,
      C_S02_AXIS_FIFO_MODE => 0,
      C_S02_AXIS_IS_ACLK_ASYNC => 0,
      C_S02_AXIS_REG_CONFIG => 0,
      C_S02_AXIS_TDATA_WIDTH => 8,
      C_S02_AXIS_TUSER_WIDTH => 1,
      C_S03_AXIS_ACLK_RATIO => 12,
      C_S03_AXIS_FIFO_DEPTH => 32,
      C_S03_AXIS_FIFO_MODE => 0,
      C_S03_AXIS_IS_ACLK_ASYNC => 0,
      C_S03_AXIS_REG_CONFIG => 0,
      C_S03_AXIS_TDATA_WIDTH => 8,
      C_S03_AXIS_TUSER_WIDTH => 1,
      C_S04_AXIS_ACLK_RATIO => 12,
      C_S04_AXIS_FIFO_DEPTH => 32,
      C_S04_AXIS_FIFO_MODE => 0,
      C_S04_AXIS_IS_ACLK_ASYNC => 0,
      C_S04_AXIS_REG_CONFIG => 0,
      C_S04_AXIS_TDATA_WIDTH => 8,
      C_S04_AXIS_TUSER_WIDTH => 1,
      C_S05_AXIS_ACLK_RATIO => 12,
      C_S05_AXIS_FIFO_DEPTH => 32,
      C_S05_AXIS_FIFO_MODE => 0,
      C_S05_AXIS_IS_ACLK_ASYNC => 0,
      C_S05_AXIS_REG_CONFIG => 0,
      C_S05_AXIS_TDATA_WIDTH => 8,
      C_S05_AXIS_TUSER_WIDTH => 1,
      C_S06_AXIS_ACLK_RATIO => 12,
      C_S06_AXIS_FIFO_DEPTH => 32,
      C_S06_AXIS_FIFO_MODE => 0,
      C_S06_AXIS_IS_ACLK_ASYNC => 0,
      C_S06_AXIS_REG_CONFIG => 0,
      C_S06_AXIS_TDATA_WIDTH => 8,
      C_S06_AXIS_TUSER_WIDTH => 1,
      C_S07_AXIS_ACLK_RATIO => 12,
      C_S07_AXIS_FIFO_DEPTH => 32,
      C_S07_AXIS_FIFO_MODE => 0,
      C_S07_AXIS_IS_ACLK_ASYNC => 0,
      C_S07_AXIS_REG_CONFIG => 0,
      C_S07_AXIS_TDATA_WIDTH => 8,
      C_S07_AXIS_TUSER_WIDTH => 1,
      C_S08_AXIS_ACLK_RATIO => 12,
      C_S08_AXIS_FIFO_DEPTH => 32,
      C_S08_AXIS_FIFO_MODE => 0,
      C_S08_AXIS_IS_ACLK_ASYNC => 0,
      C_S08_AXIS_REG_CONFIG => 0,
      C_S08_AXIS_TDATA_WIDTH => 8,
      C_S08_AXIS_TUSER_WIDTH => 1,
      C_S09_AXIS_ACLK_RATIO => 12,
      C_S09_AXIS_FIFO_DEPTH => 32,
      C_S09_AXIS_FIFO_MODE => 0,
      C_S09_AXIS_IS_ACLK_ASYNC => 0,
      C_S09_AXIS_REG_CONFIG => 0,
      C_S09_AXIS_TDATA_WIDTH => 8,
      C_S09_AXIS_TUSER_WIDTH => 1,
      C_S10_AXIS_ACLK_RATIO => 12,
      C_S10_AXIS_FIFO_DEPTH => 32,
      C_S10_AXIS_FIFO_MODE => 0,
      C_S10_AXIS_IS_ACLK_ASYNC => 0,
      C_S10_AXIS_REG_CONFIG => 0,
      C_S10_AXIS_TDATA_WIDTH => 8,
      C_S10_AXIS_TUSER_WIDTH => 1,
      C_S11_AXIS_ACLK_RATIO => 12,
      C_S11_AXIS_FIFO_DEPTH => 32,
      C_S11_AXIS_FIFO_MODE => 0,
      C_S11_AXIS_IS_ACLK_ASYNC => 0,
      C_S11_AXIS_REG_CONFIG => 0,
      C_S11_AXIS_TDATA_WIDTH => 8,
      C_S11_AXIS_TUSER_WIDTH => 1,
      C_S12_AXIS_ACLK_RATIO => 12,
      C_S12_AXIS_FIFO_DEPTH => 32,
      C_S12_AXIS_FIFO_MODE => 0,
      C_S12_AXIS_IS_ACLK_ASYNC => 0,
      C_S12_AXIS_REG_CONFIG => 0,
      C_S12_AXIS_TDATA_WIDTH => 8,
      C_S12_AXIS_TUSER_WIDTH => 1,
      C_S13_AXIS_ACLK_RATIO => 12,
      C_S13_AXIS_FIFO_DEPTH => 32,
      C_S13_AXIS_FIFO_MODE => 0,
      C_S13_AXIS_IS_ACLK_ASYNC => 0,
      C_S13_AXIS_REG_CONFIG => 0,
      C_S13_AXIS_TDATA_WIDTH => 8,
      C_S13_AXIS_TUSER_WIDTH => 1,
      C_S14_AXIS_ACLK_RATIO => 12,
      C_S14_AXIS_FIFO_DEPTH => 32,
      C_S14_AXIS_FIFO_MODE => 0,
      C_S14_AXIS_IS_ACLK_ASYNC => 0,
      C_S14_AXIS_REG_CONFIG => 0,
      C_S14_AXIS_TDATA_WIDTH => 8,
      C_S14_AXIS_TUSER_WIDTH => 1,
      C_S15_AXIS_ACLK_RATIO => 12,
      C_S15_AXIS_FIFO_DEPTH => 32,
      C_S15_AXIS_FIFO_MODE => 0,
      C_S15_AXIS_IS_ACLK_ASYNC => 0,
      C_S15_AXIS_REG_CONFIG => 0,
      C_S15_AXIS_TDATA_WIDTH => 8,
      C_S15_AXIS_TUSER_WIDTH => 1,
      C_SWITCH_ACLK_RATIO => 12,
      C_SWITCH_MAX_XFERS_PER_ARB => 1,
      C_SWITCH_MI_REG_CONFIG => 0,
      C_SWITCH_MODE => 1,
      C_SWITCH_NUM_CYCLES_TIMEOUT => 0,
      C_SWITCH_SIGNAL_SET => X"13",
      C_SWITCH_SI_REG_CONFIG => 1,
      C_SWITCH_TDATA_WIDTH => 8,
      C_SWITCH_TDEST_WIDTH => 1,
      C_SWITCH_TID_WIDTH => 1,
      C_SWITCH_TUSER_WIDTH => 1,
      C_SWITCH_USE_ACLKEN => 0
    )
    PORT MAP (
      ACLK => ACLK,
      ARESETN => ARESETN,
      ACLKEN => '0',
      S00_AXIS_ACLK => S00_AXIS_ACLK,
      S01_AXIS_ACLK => '0',
      S02_AXIS_ACLK => '0',
      S03_AXIS_ACLK => '0',
      S04_AXIS_ACLK => '0',
      S05_AXIS_ACLK => '0',
      S06_AXIS_ACLK => '0',
      S07_AXIS_ACLK => '0',
      S08_AXIS_ACLK => '0',
      S09_AXIS_ACLK => '0',
      S10_AXIS_ACLK => '0',
      S11_AXIS_ACLK => '0',
      S12_AXIS_ACLK => '0',
      S13_AXIS_ACLK => '0',
      S14_AXIS_ACLK => '0',
      S15_AXIS_ACLK => '0',
      S00_AXIS_ARESETN => S00_AXIS_ARESETN,
      S01_AXIS_ARESETN => '0',
      S02_AXIS_ARESETN => '0',
      S03_AXIS_ARESETN => '0',
      S04_AXIS_ARESETN => '0',
      S05_AXIS_ARESETN => '0',
      S06_AXIS_ARESETN => '0',
      S07_AXIS_ARESETN => '0',
      S08_AXIS_ARESETN => '0',
      S09_AXIS_ARESETN => '0',
      S10_AXIS_ARESETN => '0',
      S11_AXIS_ARESETN => '0',
      S12_AXIS_ARESETN => '0',
      S13_AXIS_ARESETN => '0',
      S14_AXIS_ARESETN => '0',
      S15_AXIS_ARESETN => '0',
      S00_AXIS_ACLKEN => '0',
      S01_AXIS_ACLKEN => '0',
      S02_AXIS_ACLKEN => '0',
      S03_AXIS_ACLKEN => '0',
      S04_AXIS_ACLKEN => '0',
      S05_AXIS_ACLKEN => '0',
      S06_AXIS_ACLKEN => '0',
      S07_AXIS_ACLKEN => '0',
      S08_AXIS_ACLKEN => '0',
      S09_AXIS_ACLKEN => '0',
      S10_AXIS_ACLKEN => '0',
      S11_AXIS_ACLKEN => '0',
      S12_AXIS_ACLKEN => '0',
      S13_AXIS_ACLKEN => '0',
      S14_AXIS_ACLKEN => '0',
      S15_AXIS_ACLKEN => '0',
      S00_AXIS_TVALID => S00_AXIS_TVALID,
      S01_AXIS_TVALID => '0',
      S02_AXIS_TVALID => '0',
      S03_AXIS_TVALID => '0',
      S04_AXIS_TVALID => '0',
      S05_AXIS_TVALID => '0',
      S06_AXIS_TVALID => '0',
      S07_AXIS_TVALID => '0',
      S08_AXIS_TVALID => '0',
      S09_AXIS_TVALID => '0',
      S10_AXIS_TVALID => '0',
      S11_AXIS_TVALID => '0',
      S12_AXIS_TVALID => '0',
      S13_AXIS_TVALID => '0',
      S14_AXIS_TVALID => '0',
      S15_AXIS_TVALID => '0',
      S00_AXIS_TREADY => S00_AXIS_TREADY,
      S00_AXIS_TDATA => S00_AXIS_TDATA,
      S01_AXIS_TDATA => (others => '0'),
      S02_AXIS_TDATA => (others => '0'),
      S03_AXIS_TDATA => (others => '0'),
      S04_AXIS_TDATA => (others => '0'),
      S05_AXIS_TDATA => (others => '0'),
      S06_AXIS_TDATA => (others => '0'),
      S07_AXIS_TDATA => (others => '0'),
      S08_AXIS_TDATA => (others => '0'),
      S09_AXIS_TDATA => (others => '0'),
      S10_AXIS_TDATA => (others => '0'),
      S11_AXIS_TDATA => (others => '0'),
      S12_AXIS_TDATA => (others => '0'),
      S13_AXIS_TDATA => (others => '0'),
      S14_AXIS_TDATA => (others => '0'),
      S15_AXIS_TDATA => (others => '0'),
      S00_AXIS_TSTRB => (others => '0'),
      S01_AXIS_TSTRB => (others => '0'),
      S02_AXIS_TSTRB => (others => '0'),
      S03_AXIS_TSTRB => (others => '0'),
      S04_AXIS_TSTRB => (others => '0'),
      S05_AXIS_TSTRB => (others => '0'),
      S06_AXIS_TSTRB => (others => '0'),
      S07_AXIS_TSTRB => (others => '0'),
      S08_AXIS_TSTRB => (others => '0'),
      S09_AXIS_TSTRB => (others => '0'),
      S10_AXIS_TSTRB => (others => '0'),
      S11_AXIS_TSTRB => (others => '0'),
      S12_AXIS_TSTRB => (others => '0'),
      S13_AXIS_TSTRB => (others => '0'),
      S14_AXIS_TSTRB => (others => '0'),
      S15_AXIS_TSTRB => (others => '0'),
      S00_AXIS_TKEEP => (others => '0'),
      S01_AXIS_TKEEP => (others => '0'),
      S02_AXIS_TKEEP => (others => '0'),
      S03_AXIS_TKEEP => (others => '0'),
      S04_AXIS_TKEEP => (others => '0'),
      S05_AXIS_TKEEP => (others => '0'),
      S06_AXIS_TKEEP => (others => '0'),
      S07_AXIS_TKEEP => (others => '0'),
      S08_AXIS_TKEEP => (others => '0'),
      S09_AXIS_TKEEP => (others => '0'),
      S10_AXIS_TKEEP => (others => '0'),
      S11_AXIS_TKEEP => (others => '0'),
      S12_AXIS_TKEEP => (others => '0'),
      S13_AXIS_TKEEP => (others => '0'),
      S14_AXIS_TKEEP => (others => '0'),
      S15_AXIS_TKEEP => (others => '0'),
      S00_AXIS_TLAST => S00_AXIS_TLAST,
      S01_AXIS_TLAST => '0',
      S02_AXIS_TLAST => '0',
      S03_AXIS_TLAST => '0',
      S04_AXIS_TLAST => '0',
      S05_AXIS_TLAST => '0',
      S06_AXIS_TLAST => '0',
      S07_AXIS_TLAST => '0',
      S08_AXIS_TLAST => '0',
      S09_AXIS_TLAST => '0',
      S10_AXIS_TLAST => '0',
      S11_AXIS_TLAST => '0',
      S12_AXIS_TLAST => '0',
      S13_AXIS_TLAST => '0',
      S14_AXIS_TLAST => '0',
      S15_AXIS_TLAST => '0',
      S00_AXIS_TID => (others => '0'),
      S01_AXIS_TID => (others => '0'),
      S02_AXIS_TID => (others => '0'),
      S03_AXIS_TID => (others => '0'),
      S04_AXIS_TID => (others => '0'),
      S05_AXIS_TID => (others => '0'),
      S06_AXIS_TID => (others => '0'),
      S07_AXIS_TID => (others => '0'),
      S08_AXIS_TID => (others => '0'),
      S09_AXIS_TID => (others => '0'),
      S10_AXIS_TID => (others => '0'),
      S11_AXIS_TID => (others => '0'),
      S12_AXIS_TID => (others => '0'),
      S13_AXIS_TID => (others => '0'),
      S14_AXIS_TID => (others => '0'),
      S15_AXIS_TID => (others => '0'),
      S00_AXIS_TDEST => (others => '0'),
      S01_AXIS_TDEST => (others => '0'),
      S02_AXIS_TDEST => (others => '0'),
      S03_AXIS_TDEST => (others => '0'),
      S04_AXIS_TDEST => (others => '0'),
      S05_AXIS_TDEST => (others => '0'),
      S06_AXIS_TDEST => (others => '0'),
      S07_AXIS_TDEST => (others => '0'),
      S08_AXIS_TDEST => (others => '0'),
      S09_AXIS_TDEST => (others => '0'),
      S10_AXIS_TDEST => (others => '0'),
      S11_AXIS_TDEST => (others => '0'),
      S12_AXIS_TDEST => (others => '0'),
      S13_AXIS_TDEST => (others => '0'),
      S14_AXIS_TDEST => (others => '0'),
      S15_AXIS_TDEST => (others => '0'),
      S00_AXIS_TUSER => (others => '0'),
      S01_AXIS_TUSER => (others => '0'),
      S02_AXIS_TUSER => (others => '0'),
      S03_AXIS_TUSER => (others => '0'),
      S04_AXIS_TUSER => (others => '0'),
      S05_AXIS_TUSER => (others => '0'),
      S06_AXIS_TUSER => (others => '0'),
      S07_AXIS_TUSER => (others => '0'),
      S08_AXIS_TUSER => (others => '0'),
      S09_AXIS_TUSER => (others => '0'),
      S10_AXIS_TUSER => (others => '0'),
      S11_AXIS_TUSER => (others => '0'),
      S12_AXIS_TUSER => (others => '0'),
      S13_AXIS_TUSER => (others => '0'),
      S14_AXIS_TUSER => (others => '0'),
      S15_AXIS_TUSER => (others => '0'),
      M00_AXIS_ACLK => M00_AXIS_ACLK,
      M01_AXIS_ACLK => '0',
      M02_AXIS_ACLK => '0',
      M03_AXIS_ACLK => '0',
      M04_AXIS_ACLK => '0',
      M05_AXIS_ACLK => '0',
      M06_AXIS_ACLK => '0',
      M07_AXIS_ACLK => '0',
      M08_AXIS_ACLK => '0',
      M09_AXIS_ACLK => '0',
      M10_AXIS_ACLK => '0',
      M11_AXIS_ACLK => '0',
      M12_AXIS_ACLK => '0',
      M13_AXIS_ACLK => '0',
      M14_AXIS_ACLK => '0',
      M15_AXIS_ACLK => '0',
      M00_AXIS_ARESETN => M00_AXIS_ARESETN,
      M01_AXIS_ARESETN => '0',
      M02_AXIS_ARESETN => '0',
      M03_AXIS_ARESETN => '0',
      M04_AXIS_ARESETN => '0',
      M05_AXIS_ARESETN => '0',
      M06_AXIS_ARESETN => '0',
      M07_AXIS_ARESETN => '0',
      M08_AXIS_ARESETN => '0',
      M09_AXIS_ARESETN => '0',
      M10_AXIS_ARESETN => '0',
      M11_AXIS_ARESETN => '0',
      M12_AXIS_ARESETN => '0',
      M13_AXIS_ARESETN => '0',
      M14_AXIS_ARESETN => '0',
      M15_AXIS_ARESETN => '0',
      M00_AXIS_ACLKEN => '0',
      M01_AXIS_ACLKEN => '0',
      M02_AXIS_ACLKEN => '0',
      M03_AXIS_ACLKEN => '0',
      M04_AXIS_ACLKEN => '0',
      M05_AXIS_ACLKEN => '0',
      M06_AXIS_ACLKEN => '0',
      M07_AXIS_ACLKEN => '0',
      M08_AXIS_ACLKEN => '0',
      M09_AXIS_ACLKEN => '0',
      M10_AXIS_ACLKEN => '0',
      M11_AXIS_ACLKEN => '0',
      M12_AXIS_ACLKEN => '0',
      M13_AXIS_ACLKEN => '0',
      M14_AXIS_ACLKEN => '0',
      M15_AXIS_ACLKEN => '0',
      M00_AXIS_TVALID => M00_AXIS_TVALID,
      M00_AXIS_TREADY => M00_AXIS_TREADY,
      M01_AXIS_TREADY => '0',
      M02_AXIS_TREADY => '0',
      M03_AXIS_TREADY => '0',
      M04_AXIS_TREADY => '0',
      M05_AXIS_TREADY => '0',
      M06_AXIS_TREADY => '0',
      M07_AXIS_TREADY => '0',
      M08_AXIS_TREADY => '0',
      M09_AXIS_TREADY => '0',
      M10_AXIS_TREADY => '0',
      M11_AXIS_TREADY => '0',
      M12_AXIS_TREADY => '0',
      M13_AXIS_TREADY => '0',
      M14_AXIS_TREADY => '0',
      M15_AXIS_TREADY => '0',
      M00_AXIS_TDATA => M00_AXIS_TDATA,
      M00_AXIS_TLAST => M00_AXIS_TLAST,
      S00_ARB_REQ_SUPPRESS => '0',
      S01_ARB_REQ_SUPPRESS => '0',
      S02_ARB_REQ_SUPPRESS => '0',
      S03_ARB_REQ_SUPPRESS => '0',
      S04_ARB_REQ_SUPPRESS => '0',
      S05_ARB_REQ_SUPPRESS => '0',
      S06_ARB_REQ_SUPPRESS => '0',
      S07_ARB_REQ_SUPPRESS => '0',
      S08_ARB_REQ_SUPPRESS => '0',
      S09_ARB_REQ_SUPPRESS => '0',
      S10_ARB_REQ_SUPPRESS => '0',
      S11_ARB_REQ_SUPPRESS => '0',
      S12_ARB_REQ_SUPPRESS => '0',
      S13_ARB_REQ_SUPPRESS => '0',
      S14_ARB_REQ_SUPPRESS => '0',
      S15_ARB_REQ_SUPPRESS => '0'
    );

END spartan6;
