library ieee;
use ieee.STD_LOGIC_1164.ALL;

use ieee.NUMERIC_STD.ALL;

entity process_trigger_TB is
end entity;

architecture test_bench of process_trigger_TB is


  
signal clk
    signal rst
    signal data_input
    signal scaler_count
    signal scaler_count_pixel
    signal new_hit


end architecture;     
